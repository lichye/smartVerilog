//# 62 inputs
//# 152 outputs
//# 638 D-type flipflops
//# 5378 inverters
//# 2573 gates (1114 ANDs + 849 NANDs + 512 ORs + 98 NORs)



module dff (CK,Q,D);
input CK,D;
output Q;
  wire NM,NCK;
  reg NQ,M; // trireg -> reg
  assign M = D ? NCK : 1'bz; //nmos N7 (M,D,NCK);
  assign NQ = NM ? CK : 1'bz; //nmos N9 (NQ,NM,CK);
  not P3 (NM,M);
  not P5 (Q,NQ);
  not P1 (NCK,CK);

endmodule



module s13207(GND,VDD,CK,g1,g10,g1000,g1006,g1008,g1015,g1016,g1017,g1080,g11,
  g1193,
  g1194,g1195,g1196,g1197,g1198,g1201,g1202,g1203,g1205,g1206,g1234,g1246,
  g1553,g1554,g1724,g1783,g1798,g1804,g1810,g1817,g1824,g1829,g1870,g1871,
  g1894,g1911,g1944,g206,g21,g22,g23,g24,g25,g26,g2662,g27,g28,g2844,g2888,g29,
  g291,g30,g3077,g3096,g31,g3130,g3159,g3191,g32,g37,g372,g3829,g3854,g3856,
  g3857,g3859,g3860,g41,g42,g4267,g43,g4316,g4370,g4371,g4372,g4373,g44,g45,
  g453,g4655,g4657,g4660,g4661,g4663,g4664,g49,g5143,g5164,g534,g5571,g5669,
  g5678,g5682,g5684,g5687,g5729,g594,g6207,g6212,g6223,g6236,g6269,g6288,g6289,
  g6290,g6291,g6292,g6293,g6294,g6295,g6296,g6297,g6298,g6299,g6300,g6301,
  g6302,g6303,g6304,g6305,g6306,g6307,g6308,g633,g634,g635,g6376,g6425,g645,
  g647,g648,g6648,g6653,g6675,g6849,g6850,g6895,g690,g6909,g694,g698,g702,
  g7048,g7063,g7103,g722,g723,g7283,g7284,g7285,g7286,g7287,g7288,g7289,g7290,
  g7291,g7292,g7293,g7294,g7295,g7298,g7423,g7424,g7425,g7474,g7504,g7505,
  g7506,g7507,g7508,g751,g7514,g752,g753,g754,g755,g756,g757,g7729,g7730,g7731,
  g7732,g7763,g781,g785,g786,g795,g8216,g8217,g8218,g8219,g8234,g8661,g8663,
  g8872,g8958,g9,g9128,g9132,g9204,g9280,g929,g9297,g9299,g9305,g9308,g9310,
  g9312,g9314,g9378,g941,g955,g962);
input GND,VDD,CK,g43,g49,g633,g634,g635,g645,g647,g648,g690,g694,g698,g702,
  g722,g723,g751,
  g752,g753,g754,g755,g756,g757,g781,g941,g962,g1000,g1008,g1016,g1080,g1234,
  g1553,g1554,g786,g1206,g929,g955,g795,g1194,g1198,g1202,g24,g1203,g1196,g29,
  g22,g28,g10,g23,g37,g26,g1,g27,g42,g11,g32,g41,g31,g45,g9,g44,g21,g30,g25;
output g206,g291,g372,g453,g534,g594,g785,g1006,g1015,g1017,g1246,g1724,g1783,
  g1798,g1804,g1810,g1817,g1824,g1829,g1870,g1871,g1894,g1911,g1944,g2662,
  g2844,g2888,g3077,g3096,g3130,g3159,g3191,g3829,g3859,g3860,g4267,g4316,
  g4370,g4371,g4372,g4373,g4655,g4657,g4660,g4661,g4663,g4664,g5143,g5164,
  g5571,g5669,g5678,g5682,g5684,g5687,g5729,g6207,g6212,g6223,g6236,g6269,
  g6425,g6648,g6653,g6675,g6849,g6850,g6895,g6909,g7048,g7063,g7103,g7283,
  g7284,g7285,g7286,g7287,g7288,g7289,g7290,g7291,g7292,g7293,g7294,g7295,
  g7298,g7423,g7424,g7425,g7474,g7504,g7505,g7506,g7507,g7508,g7514,g7729,
  g7730,g7731,g7732,g8216,g8217,g8218,g8219,g8234,g8661,g8663,g8872,g8958,
  g9128,g9132,g9204,g9280,g9297,g9299,g9305,g9308,g9310,g9312,g9314,g9378,
  g7763,g1205,g3856,g3857,g3854,g1193,g1197,g1201,g6294,g6376,g1195,g6300,
  g6292,g6298,g6291,g6293,g6304,g6296,g6289,g6297,g6306,g6290,g6303,g6305,
  g6302,g6308,g6288,g6307,g6299,g6301,g6295;

  wire g397,g4635,g1271,g5176,g312,g4618,g273,g4611,g452,g449,g948,g8664,g629,
    g6827,g207,g5733,g1541,g7778,g1153,g6856,g940,g5735,g976,g8864,g498,g9111,
    g314,g4620,g1092,g7520,g454,g4639,g196,g5731,g535,g3844,g292,g4613,g772,
    g6846,g1375,g6869,g689,g6371,g183,g6309,g359,g6336,g1384,g6881,g1339,g6865,
    g20,g6386,g1424,g3862,g767,g6841,g393,g4631,g1077,g7767,g1231,g1236,g294,
    g4615,g1477,g9036,g4,g9372,g608,g6806,g1204,g465,g6352,g774,g6848,g921,
    g916,g1304,g1312,g243,g6318,g1499,g7772,g80,g6778,g1444,g5185,g1269,g5740,
    g600,g6807,g423,g9105,g771,g6845,g803,g7757,g843,g2647,g315,g4621,g455,
    g4640,g906,g901,g622,g6821,g891,g3855,g1014,g1012,g984,g9133,g117,g5153,
    g137,g5150,g527,g9110,g1513,g1524,g278,g6323,g1378,g6880,g718,g7753,g598,
    g6797,g1182,g1160,g1288,g7527,g1382,g6888,g179,g5159,g624,g6831,g48,g9362,
    g362,g9093,g878,g890,g270,g9092,g763,g6836,g710,g7751,g730,g7754,g295,
    g4616,g1037,g7519,g1102,g6855,g483,g6356,g775,g7759,g621,g6819,g1364,g6878,
    g1454,g5187,g1296,g7304,g5,g9373,g1532,g7781,g587,g3852,g741,g9386,g13,
    g7308,g606,g6804,g6851,g52,g6781,g646,g4652,g1412,g5745,g327,g6332,g1189,
    g6392,g1389,g4658,g1029,g2654,g1371,g6868,g1429,g2671,g398,g4636,g985,
    g7515,g354,g4624,g619,g6817,g113,g5148,g133,g5149,g180,g5158,g1138,g7524,
    g1309,g1308,g889,g7101,g390,g6341,g625,g6823,g417,g9103,g681,g7748,g437,
    g6348,g351,g9100,g1200,g109,g6785,g1049,g8673,g1098,g6854,g200,g199,g240,
    g6317,g479,g4649,g126,g6789,g596,g6795,g1268,g5175,g222,g6313,g420,g9104,
    g3,g9360,g58,g7734,g172,g1270,g387,g6340,g840,g2648,g365,g9094,g1486,g8226,
    g1504,g7773,g1185,g1155,g1385,g6883,g583,g3851,g822,g7512,g1025,g8871,g969,
    g966,g768,g6842,g174,g7737,g685,g7749,g1087,g6853,g355,g4625,g911,g1226,
    g6859,g99,g6783,g1045,g8224,g1173,g7526,g1373,g6871,g186,g3830,g760,g6833,
    g959,g5169,g1369,g6875,g1007,g8867,g1459,g3863,g758,g6840,g480,g6355,g396,
    g4634,g612,g6811,g38,g5746,g632,g6830,g1415,g5180,g1227,g7108,g246,g6319,
    g3840,g517,g4651,g118,g6787,g138,g6792,g16,g1404,g284,g9086,g142,g6793,
    g219,g6312,g426,g9106,g1388,g6882,g806,g7510,g846,g2646,g1428,g2672,g579,
    g3850,g1030,g7518,g614,g6812,g1430,g4666,g1247,g6380,g669,g7745,g110,g130,
    g6790,g225,g6314,g281,g9085,g819,g7761,g6385,g611,g6810,g631,g6829,g1217,
    g6377,g104,g6784,g1365,g6867,g825,g7513,g1333,g6863,g474,g4644,g1396,g4662,
    g141,g5151,g1509,g7774,g766,g6839,g1018,g8869,g588,g9031,g1467,g8875,g317,
    g4623,g457,g4642,g486,g6357,g471,g6354,g1381,g6887,g513,g9116,g1397,g6389,
    g533,g530,g1021,g8870,g1421,g5179,g952,g8668,g1263,g5737,g580,g6368,g615,
    g6813,g1257,g5738,g46,g8955,g402,g6343,g998,g1005,g1041,g7765,g297,g6324,
    g954,g8670,g105,g145,g5152,g212,g4601,g1368,g6874,g232,g4606,g990,g7516,
    g475,g4645,g33,g5184,g951,g8667,g799,g7756,g812,g7758,g567,g6367,g313,
    g4619,g333,g6334,g168,g7742,g214,g4603,g234,g4608,g652,g1126,g8674,g1400,
    g6390,g1326,g7306,g92,g6794,g309,g6328,g211,g4600,g834,g2650,g231,g4605,
    g557,g6366,g1383,g6889,g1220,g6378,g158,g7740,g627,g6825,g661,g7743,g77,
    g6777,g831,g2651,g1327,g7307,g293,g4614,g1146,g1612,g89,g150,g7738,g773,
    g6847,g859,g8221,g1240,g1235,g518,g6361,g1472,g8960,g1443,g4667,g436,g4638,
    g405,g6344,g1034,g8957,g1147,g374,g4627,g98,g5146,g563,g9029,g510,g9115,
    g3842,g215,g4604,g235,g4609,g1013,g6,g9374,g55,g7733,g1317,g5743,g504,
    g9113,g665,g7744,g544,g6365,g371,g368,g62,g7509,g792,g5162,g468,g6353,g815,
    g7760,g1460,g4668,g553,g9028,g623,g6822,g501,g9112,g1190,g8677,g1390,g4659,
    g74,g6776,g1156,g1081,g318,g6329,g458,g4643,g342,g9097,g1250,g7111,g1163,
    g2655,g1363,g6877,g1432,g5183,g1053,g8873,g252,g6321,g330,g6333,g264,g9090,
    g1157,g1357,g8675,g375,g4628,g68,g6774,g852,g2644,g261,g9089,g516,g4650,
    g536,g6363,g979,g7104,g778,g7296,g3832,g1292,g7302,g290,g287,g1084,g7106,
    g1439,g5182,g770,g6844,g1276,g6384,g7102,g1004,g7105,g1403,g93,g5145,g2,
    g9361,g3836,g560,g6370,g1224,g6857,g1320,g7114,g617,g6815,g316,g4622,g336,
    g9095,g933,g5166,g456,g4641,g345,g9098,g628,g6826,g8,g9376,g887,g7099,g789,
    g7297,g173,g7736,g550,g9027,g255,g9087,g949,g8665,g1244,g2659,g620,g6818,
    g1435,g5181,g477,g4647,g926,g3838,g855,g8220,g1214,g5736,g1110,g7299,g1310,
    g296,g4617,g972,g2653,g1402,g6391,g896,g613,g6820,g566,g3848,g1394,g6388,
    g1489,g7770,g883,g47,g9389,g971,g5171,g609,g6808,g103,g5157,g1254,g6381,
    g556,g3847,g1409,g5178,g626,g6824,g1229,g7110,g782,g5734,g237,g6316,g942,
    g2652,g228,g6315,g706,g7750,g746,g8956,g1462,g8678,g963,g7764,g129,g5156,
    g837,g2649,g599,g6798,g1192,g1191,g828,g7762,g1392,g6387,g492,g6359,g95,
    g94,g944,g6372,g195,g3831,g1431,g2673,g1252,g2661,g356,g6335,g953,g8669,
    g1176,g5172,g1376,g6890,g1405,g5744,g1225,g6858,g1073,g9145,g1324,g7118,
    g1069,g9134,g443,g9101,g1377,g6891,g377,g4630,g618,g6816,g602,g6800,g213,
    g4602,g233,g4607,g1199,g6375,g1399,g3861,g83,g6779,g888,g7100,g573,g9033,
    g399,g6342,g1245,g507,g9114,g547,g9026,g108,g5147,g610,g6809,g630,g6828,
    g1207,g5173,g249,g6320,g65,g4598,g936,g5168,g478,g4648,g604,g6802,g945,
    g5170,g1114,g7521,g100,g429,g9107,g809,g7511,g849,g2645,g1408,g5177,g1336,
    g6864,g601,g6799,g122,g6788,g1065,g9117,g1122,g8225,g1228,g7109,g495,g6360,
    g1322,g7116,g1230,g7300,g1033,g9034,g267,g9091,g6374,g1395,g1393,g373,
    g4626,g274,g4612,g1266,g5739,g714,g7752,g734,g7755,g1142,g8874,g1342,g7119,
    g769,g6843,g6852,g1481,g7769,g1097,g543,g3846,g1154,g1354,g7768,g489,g6358,
    g874,g4654,g121,g5154,g591,g9032,g616,g6814,g1267,g4656,g1311,g605,g6803,
    g182,g5161,g1401,g950,g8666,g1329,g2663,g408,g6345,g871,g5167,g759,g6832,
    g146,g7735,g202,g5732,g440,g6349,g476,g4646,g184,g6310,g1149,g7525,g1398,
    g210,g3834,g394,g4632,g86,g6780,g570,g9030,g275,g6322,g303,g6326,g125,
    g5155,g181,g5160,g6393,g595,g576,g1319,g7113,g863,g8222,g1211,g5174,g8223,
    g1186,g1386,g6884,g875,g5165,g1170,g1370,g6876,g201,g1325,g7305,g1280,
    g7112,g1106,g7107,g1061,g9035,g1387,g6885,g762,g6835,g1461,g4669,g378,
    g6337,g1514,g7775,g1345,g7528,g6373,g1391,g185,g4599,g1307,g3858,g1159,
    g1223,g6379,g446,g9102,g1416,g4665,g395,g4633,g764,g6837,g1251,g6860,g216,
    g6311,g236,g4610,g205,g3835,g540,g6364,g3849,g1537,g7777,g727,g8228,g999,
    g8865,g761,g6834,g1272,g6383,g1243,g2660,g1328,g7309,g1130,g7522,g1330,
    g6862,g114,g6786,g134,g6791,g1166,g1167,g524,g9109,g1366,g6866,g348,g9099,
    g1148,g1348,g7529,g1260,g6382,g7,g9375,g258,g9088,g521,g6362,g300,g6325,
    g765,g6838,g1118,g7766,g1318,g6861,g1367,g6873,g677,g7747,g376,g4629,g1057,
    g8959,g973,g8672,g2664,g1549,g7780,g1321,g7115,g1253,g5741,g1519,g8227,
    g584,g6369,g539,g3845,g324,g6331,g432,g9108,g1158,g321,g6330,g414,g6347,
    g1374,g6872,g6782,g1284,g7301,g1545,g7779,g1380,g6886,g673,g7746,g607,
    g6805,g306,g6327,g943,g8671,g162,g7741,g411,g6346,g866,g5163,g1300,g7303,
    g384,g6339,g339,g9096,g459,g6350,g1323,g7117,g381,g6338,g1528,g7776,g1351,
    g7530,g597,g6796,g1372,g6870,g154,g7739,g435,g4637,g970,g1134,g7523,g995,
    g7517,g190,g1313,g5742,g603,g6801,g1494,g7771,g462,g6351,g1360,g8676,g1450,
    g5186,g187,g5730,g1179,g1379,g6879,g12,g8662,g71,g6775,g1658,g1777,I9325,
    g4242,I7758,g2605,g5652,I10135,I13502,g7135,I12558,g3880,g2965,I12382,
    I15824,g9157,g5843,g5367,I6112,g7189,I13109,g8970,I15414,I6267,g6062,
    I10675,I16126,g9354,I10519,g5242,I15181,g8734,I11443,g6038,I12436,g6635,
    g5662,g2547,I6371,I7365,g3061,I10154,g5109,g1611,I11278,g5780,g7171,g7071,
    I14154,g7558,I12274,g6672,I14451,g5834,I10525,g5971,I10587,g3978,g3160,
    I6676,g1603,g3612,I7082,I8520,g3652,g2892,g2266,I13469,g7123,I12346,g6737,
    I9636,g4802,I14637,g8012,I12235,g1799,I5657,g3935,I7602,I5933,g9207,g9197,
    I13039,g6961,I15426,g8895,g5598,g4938,g1674,g7281,I13277,g3982,g3192,I8913,
    I15190,g8685,g2945,g2364,g5121,I9515,g3128,I6839,g3629,g2424,I13323,g5670,
    I10157,I11815,g6169,I12397,I6849,I15654,g8789,g8564,g3542,I12292,g6657,
    I11221,g2709,g1747,I11677,g6076,I11503,I8859,I8829,g4029,I15546,g9007,
    g1680,I5515,I15211,g8808,g2340,I12409,g6398,I8880,I14106,g7138,I12996,
    I6703,g1983,g5938,g5412,g8771,g2478,g5813,I10472,g7338,I13432,g2907,g2289,
    g1744,g9215,I15921,I12915,I12433,I12635,g6509,I13359,g1802,I10439,g5214,
    g2959,g1926,I14728,g8152,I8733,g3996,I14439,g8063,g2517,I6348,g4010,g3097,
    I7662,g3642,I9446,g3926,I8974,g3871,I10277,g5519,I9929,I15732,g1558,I5435,
    I7290,g2936,g2876,g2231,I16058,I11884,g6091,I9145,g4264,I6468,g1917,g5606,
    g4748,I8796,g3934,I14148,I14349,g7588,I11410,g5845,I12164,g5847,g695,I5392,
    g6708,g6250,I13410,g7274,I15625,g9000,g6520,I11704,g1901,I5781,g6219,
    I10998,g6640,I11908,I8980,g4535,g3902,I7495,I12891,g6950,I11479,g6201,
    I11666,g5772,I10190,g2915,I6643,I13666,g7238,g6252,g5418,I12307,I8357,
    g7049,I12813,g3512,g1616,I13478,g7126,g5586,g6958,I12675,I15943,g9214,
    I8769,I6716,g1721,I11455,I8916,I5981,I8177,g2810,I7847,g3798,I16055,g9291,
    g9336,I16084,g2310,I6087,g7715,I14022,g1600,g1574,g1864,g4566,g2902,I11556,
    g6065,g7098,g6525,I5997,I12358,g7498,I13672,I6460,I12108,g5939,g6765,g3529,
    g2323,I15391,I6198,g4693,I13580,g7208,g4134,g3676,g3649,I14139,g7548,I9416,
    g4273,I12283,g6692,g8482,g8094,g5525,g4934,I7356,g5645,I5353,g3833,g2402,
    I7950,g2774,g2824,g1688,g1580,g2236,I5969,g7584,I13897,g4555,g2894,g9065,
    I15589,I9642,g4788,g7539,I13797,I15411,g8897,I15527,g9020,I10415,g5397,
    I13084,g9322,g9313,g3964,g4792,I9111,g9230,I15950,g6225,I11014,I8781,g3932,
    I8898,g4089,g6073,g5384,g2877,g2232,I12259,g1736,I5577,I12091,g5988,I8778,
    g5607,I15513,g7162,I13060,g7268,I13244,g7019,I12771,I11740,g6136,g7362,
    I9600,I13740,g7364,I9654,I15894,g9195,I11299,I7723,g3052,g4113,g6069,
    I10690,g2556,g1889,I7101,I5901,g2222,I5939,I13676,g7256,I15678,I8291,
    I13373,g7270,g2928,g2326,g4202,I14783,I7605,g2752,I15714,g9077,g5587,g2930,
    g2328,I15315,g8738,I11800,g6164,I5754,g4908,g4088,I11458,g6206,g5639,g5311,
    g2899,g2272,I15871,g4094,I7905,I11936,g5918,g3872,g2954,I15202,g8797,I7132,
    g4567,g2903,g7728,I14055,g7486,I13646,g3843,I7332,g3989,g3131,I6186,I14061,
    I9612,g4776,I10608,g5701,I9648,g8762,g8585,I13692,I15978,g9235,I14115,
    g7563,g7185,I13099,I9081,I7041,g2401,I12418,I9935,g4812,g4593,g2939,I11964,
    g3549,g2404,I7305,g3971,I7688,g7070,g6562,g2295,I14052,g7494,g2237,I5972,
    g7470,g7253,I15741,g9083,g8657,I14763,I12214,I13550,I9666,I6574,I8215,
    g3577,g6898,I12567,g1838,g5591,g4841,g6900,I12571,I14445,I8886,g4308,g5832,
    I14813,g8640,g1795,I5649,I12262,g1737,g2394,I6270,g9248,g1809,I10973,g5726,
    I14798,g8605,g6245,g5690,g4360,I8333,I7368,g3018,g9255,I15985,g9081,I15635,
    I12948,g6919,I13909,g7339,I15735,g9078,g4521,g2866,I14184,g7726,g1672,
    I14674,g7788,g8464,g8039,I11200,I12702,g6497,g2557,g4050,g3080,I8838,
    I12757,g6577,I15681,g2966,g1856,g5794,I10421,I5889,g1643,I11569,g6279,
    g7131,g6976,I11359,g2471,I6309,g7006,I12748,g7331,I13413,I15196,g8778,
    I6636,g1704,I14732,g8155,g2242,I10962,g3909,I7520,I11747,g6123,I12564,
    g6720,g8563,I14662,g2948,g2366,I11242,g6183,I14169,I12328,I12903,g3519,
    g2185,I10761,g5302,I13347,I7856,g3805,I7734,g2595,g2955,g7487,I13649,g5628,
    g1742,g6088,I10708,I12427,g5515,g4923,g6764,g6488,I11652,I8889,g4777,I9084,
    I10400,g5201,g5100,I9484,I9512,g3985,I13807,g7320,I11974,g5956,I12062,
    I14400,g7677,g2350,I6166,I15726,I14136,g9218,I15930,I9823,g5138,I16052,
    g2038,g4882,g4069,I14214,g7576,I12933,g7018,I9366,g4350,g7226,g6937,I11230,
    g6140,I11293,g5824,I10207,g5075,I13293,g7159,I12508,g6593,I11638,I12529,
    I6446,g1812,I8748,I5356,I14005,g7434,g7045,g6490,I11416,g5829,I10538,g5255,
    I6003,I9148,g4354,I13416,g7165,I5795,g9129,I15765,g2769,g7173,g6980,g9329,
    g9317,I11269,g7091,g7491,I13653,I12481,I7383,g2918,g3341,I6936,I5839,g6650,
    g6213,g7169,I13075,I13281,g1572,I15379,I6695,g2246,g4541,g2883,g7059,g6538,
    g7920,I14282,g7578,I13879,g6008,I11835,g6181,g3691,I7195,g5621,g7459,
    I13617,g9221,I15937,I12205,I9463,g3942,g7718,I14031,I14172,g4153,I8024,
    g4680,I8945,g3650,I10773,g4353,g3665,I11586,g6256,I12912,I11335,I14100,
    g7580,I6223,g8038,g7694,g6768,I12173,g4306,g7582,I13891,g6594,I11796,g1961,
    g3879,g2963,I9129,g7261,I13225,I14683,g7825,g3962,I9579,g7793,I14234,g3158,
    I6853,g3659,g2293,I12289,g5648,I6416,g1794,g3506,g1781,g7015,I12763,I12592,
    g4558,g2897,g9068,I15598,I7126,g2494,I5926,I7400,g3075,g3968,I7326,g2940,
    I6115,I6251,g2921,g2312,I10684,I12532,g6122,I10752,I10882,g5600,g6228,
    I11021,g3587,g1964,I11275,g5768,I9457,g3940,g8918,I15340,I16180,g9387,
    g6230,I11025,g7246,I13196,g8967,I15405,I13746,g7311,I13493,g7132,I9393,
    g4266,g4511,g2841,I15660,g9062,g2895,g2268,g6033,g2837,g1780,g7721,g7344,
    g5839,I10532,I9834,g4782,g4092,I7899,I13035,g6964,I7712,I12731,g6579,
    I11806,g6275,I8715,g3465,g4574,g3466,g6096,g5317,g6496,I11662,g1679,I5512,
    I8097,g3237,g5278,I9794,I12406,g7502,I13682,I15550,g9008,g9198,g9187,g3545,
    g2344,I8354,g738,I5404,g6195,I10940,g5618,g5015,g6137,I10776,I12544,I9555,
    g1831,I11338,g3591,g1789,I7299,g4580,g2919,g9241,I15971,I7588,g2584,g3853,
    I7362,I14725,g8145,g7188,I13106,I10592,g2842,g2209,I9938,g4878,I10758,
    g1805,I5667,g1916,g5693,I10204,g7216,I13152,g1749,g2298,I6072,I14082,
    I12448,g2392,I13193,g7007,g2485,I11362,g5821,g7028,I13362,g7265,g3931,
    I7592,I8218,g3002,I15773,g9126,I6629,g2052,I8784,g7247,I13199,I5654,I6130,
    g4076,I7859,g9319,g9309,g5489,g2941,g2349,I9606,g4687,I11353,g3905,I13475,
    g7125,I14848,g8625,g6255,I11066,I12316,I10804,g5526,I6800,g2016,I9687,
    g4822,g3630,I7095,g6481,I11641,I14804,I14094,I8868,g5113,I9499,I12008,
    g6097,g5345,I11437,g5801,I15839,g9168,g2520,g9209,g2640,g1584,g9211,I15909,
    I11389,g4285,I8233,I8727,g3944,g9186,I15836,I5679,g4500,g2832,I16176,g6960,
    I12681,I15965,g9219,I7944,g3774,g1579,g703,g1869,g4960,I13356,I11347,g5761,
    g2958,g2377,g7224,I15492,I5831,g2376,I6226,g5494,I9918,g3750,g2177,I9570,
    g4696,I10406,g5203,I9341,g4251,g5719,g1752,I14406,g7681,g3973,I9525,g4413,
    I11781,g6284,I12768,g6718,I15619,g8998,g9370,I16138,I9645,g4900,I15557,
    g9010,g2829,g1785,g9125,I15753,g4024,I11236,g6148,g2286,I6042,I12220,
    I14145,g7066,I12839,I10500,g5234,I16168,g9381,g7589,I13912,I6090,g2911,
    g2292,g4795,I9116,I8932,g4096,I5422,g7466,I13622,g4809,g6267,I11086,I11263,
    g3969,I14049,g7493,I16006,I11821,g6170,I12881,g6478,g1786,g7365,I13509,
    I12810,I7347,g2985,I15641,g2270,I6015,g4477,I8517,g7448,I13605,I13063,
    g6973,g7711,I14012,g4523,g2868,g6676,I11984,I11790,g6282,I11206,I13264,
    g7061,I6148,g7055,g6517,I14436,I8844,g3666,g2134,I9158,g4256,I13137,g7027,
    g2225,I5948,g6129,g7455,I13613,I11314,g6761,I12154,g2073,g7133,I12983,
    I7697,I15708,g7333,I13419,I13873,g7342,g9306,I16036,I12355,g1770,I14193,
    g5521,g4929,I15388,I12361,I8817,g3648,g3875,g2324,g3530,g4232,g7196,I13122,
    g4742,I9064,g9061,I15577,I15601,g8992,g4104,I7925,I10605,g5440,I11422,
    g5842,g6592,g3655,g1844,I15187,g8682,I14273,g7631,I11209,g6139,I13422,
    g7586,I13209,g6912,g2540,I9615,g4739,g6221,I11004,I12003,g6202,g8765,g8524,
    g7538,I13794,I13834,I6463,g1769,I10463,g5220,g9324,I14211,I15495,g5724,
    g4969,I6229,I14463,g8072,I12779,g6740,I9663,g6703,I12041,I13707,g4926,
    g9212,g9200,g9189,g5627,g7614,g3884,I7417,g3839,I7320,g2287,I6045,g7067,
    g6658,g8974,I7317,g2893,g5658,I15791,g9140,g7418,I13533,g6624,I11864,g7467,
    g7236,g6953,g6745,I6118,I14795,g8604,I14454,g5835,I10528,I13302,I8754,
    g6068,I10687,g1888,I6872,g4044,g6468,I11622,I12945,I9591,g4710,g4444,I8452,
    g1787,I6652,I11607,g5767,I6057,I12826,g6441,I12999,g7029,I11320,g5797,
    I15666,g9070,I13320,g7139,I6457,g1886,I13659,g1675,g6677,I11987,g7058,
    I13274,g6917,I7775,g3705,g5611,g8324,I14573,g4572,g2909,I7922,g3462,g2898,
    g2271,I15478,g8910,g2900,g2273,I12469,I12672,g6473,I7581,I15711,g4543,
    g2885,g5208,I11464,g5799,I10436,I13565,g7181,g4778,I6834,g9307,g9300,g2510,
    g639,I5374,g2245,g6149,I10810,g3988,I6686,I11374,g5674,g5042,g8177,I14410,
    g3693,I11034,g5644,g9223,I14163,g7533,g2291,g7438,I12415,I15580,g8985,
    I12331,g6704,g5541,g4814,g3548,g1684,g1745,g6198,g5335,g1639,I11515,I10541,
    g5256,I6121,g7263,I13231,g2207,I5920,I9585,g5680,g5101,I12897,g6962,g6569,
    I12961,g6921,g4301,I9630,g4867,I14789,g8544,g2259,g4014,I7769,I7079,g2532,
    I12505,g6612,g9315,I16061,g1808,g4885,g4070,I13635,g7243,I10289,g8199,
    I14424,g9047,I15543,g5802,I10445,I8895,g2923,I6657,I12717,g6543,g1707,
    I14325,g7713,I10829,g5224,g8781,I10535,g5254,I5389,I5706,g8898,I15308,
    g4903,g4084,g7562,I13858,I15178,g8753,I10946,g5563,I15003,g6524,I11710,
    I14828,g8639,g6644,g6208,g8510,I14643,I13164,g7086,I5371,g7723,I14042,
    I14121,g7587,g2215,I15953,I11284,g2886,g2240,g3908,I7517,I13335,g2843,
    g7336,g9057,g4036,g6152,I10815,g6258,g5427,I11383,I12325,g1575,g1865,I8483,
    g3641,I12472,g3567,g2407,I15417,g8893,g1715,I5559,g2314,I6099,I9440,I14291,
    g7680,g6632,g4335,I9123,g4455,I15334,g8800,I14124,g2870,g5492,g4919,I12148,
    g4382,I8373,g1833,g5128,I13537,g7152,g5574,I8790,g4020,g6211,g2825,I6553,
    I6434,g6186,I10919,I11485,I12646,g6493,g7585,I13900,g9017,I15475,g4931,
    I15762,g9039,I12343,g6731,g4805,I9136,g6975,I12712,g4916,g4022,I7785,g3965,
    I7676,I5963,g6599,I11809,g1896,g7441,I15423,g8894,g6026,I9528,g4006,g6426,
    I11559,I6860,g3264,I6900,I7053,g2452,I6341,I10506,g5236,g5580,g9234,I15956,
    I10028,g4825,g6614,I11838,I14028,g7501,g3933,I8904,g4126,g9330,I11302,
    I12334,g3521,g4560,I8446,g3014,g3050,I6788,I7115,g9201,g9006,I10265,g2943,
    g2362,g6984,I12725,g7168,I13072,g6939,I7731,g6287,I12412,g6404,I8841,g3979,
    g5623,I14187,g6083,I10702,g6649,I5957,g2887,g2241,g4873,I9217,I8811,g7531,
    I13773,g4095,I7908,g5076,I8763,g3947,g4037,g2845,g6483,I11645,I12229,g6659,
    I9884,g4868,g2934,g5476,g4907,g4653,I8874,I6358,g4102,I7919,g6636,I11900,
    I15568,g8981,I15747,g9042,I5865,g9213,I15915,g6106,I9651,g4579,I10649,
    g5657,I12011,I11245,I5715,I13695,g5871,I10558,g3878,g2962,g8008,g7559,
    g4719,I9021,I12241,I14073,I6587,g1708,g3777,g2170,g7411,g7202,I9372,I10491,
    g5231,I15814,g9154,I7308,I16116,g9350,I11488,I11522,g2096,I9618,I12582,
    g5285,g6461,g8768,I13663,g7235,g3882,g2970,g2496,I7626,g3632,g4917,I15974,
    I6615,g6756,I12141,g8972,I15420,I10770,g5441,I12310,g6723,g1897,g6622,
    I11858,I13628,I8757,g3921,g6027,g7992,g7557,g4265,g3611,g6427,I11562,g2137,
    g2891,g2265,I9678,I15638,g8978,g9366,g2913,g2307,I12379,g5139,I9543,I9837,
    g6904,I12958,g6920,g9056,I15562,g8065,I14338,I8315,g6446,I11591,g3981,
    I7706,g5024,I9360,g6514,I11696,I6239,g3674,I7164,g2807,g1782,I5362,g3841,
    I11326,g5819,g4892,g5795,I10424,I10268,g8917,g6403,I13326,g7176,g5809,
    I10460,I5419,I9804,I10262,g5551,I7683,g2573,g3997,I12742,g6590,I12394,
    I15510,g8969,I11040,g5299,I11948,g5897,g6763,I12158,I7778,g3019,I16142,
    I11500,I5410,g4296,g3790,g3238,I6894,I9621,g4732,g5477,g9260,I15990,g5523,
    g6469,I10719,g5559,g6637,I11903,g5643,I10128,I15014,g8607,g1801,g4553,
    g9063,I15583,I11248,I15586,g8987,I15007,g8627,g4303,I14718,g8068,g3802,
    g1832,g7688,g7406,I11404,I11008,g2481,I6317,g8913,I15329,g1748,g2692,g1671,
    g4012,I7765,I12445,I10283,I9974,g5099,g2497,I12690,g6467,g2354,I6178,
    I16165,g9377,g2960,g2381,g4706,I9005,I9567,I7526,I5897,g8179,I10247,g5266,
    g3901,I7492,g7000,g7137,I15720,g9053,g9318,g9304,g9367,I16129,I11933,
    I12968,I8935,g4005,I5425,I7800,g6251,I11060,I11272,I12304,g6642,I11912,
    I11851,g6277,g3511,g5754,g5403,I15565,g9261,I14151,I14388,g7605,I7850,
    g2795,g9193,g9181,g3092,I6826,I14777,g8511,g3492,I6970,g4281,g2562,I12493,
    g5613,I14251,g7541,g3574,g1771,g3864,g8342,g8856,g2267,I6006,I6093,g6654,
    I11942,g5444,g5074,g5269,I9791,I7702,g3062,I15684,g9067,g8481,I12128,g1578,
    g699,g1868,I5747,g4257,g3761,I10032,g1718,I5562,I14208,I12511,g4684,I8949,
    I9050,g3881,I11452,g6071,g6595,I8832,I5682,I5766,I11047,g5653,I13574,g7205,
    g2329,I6440,g1806,g7023,g9121,g4963,g4328,g2761,g1820,I5801,g9321,g9311,
    I15394,I13544,g1582,I11311,g5760,g7359,I13311,g2828,g1980,I12298,g6697,
    I6323,g7546,g1793,I7561,I10766,g2727,g4808,g6978,I11832,g7161,I13057,I5416,
    g5144,g6243,I11050,g7361,I13499,I15193,g8774,I13051,g6967,g6969,g2746,
    I12737,g6460,g2221,I5936,g3076,g7127,g6974,g8783,g7327,I13403,I12232,g6662,
    g1664,I6151,g2703,I14433,I8823,g5014,I9344,g6130,g7146,g6998,g6542,I11718,
    I11317,g7346,I13454,g7633,I13962,I5565,I11350,g5763,g2953,I7970,g3557,
    I13350,g7223,g8901,g2932,I9271,g4263,g3651,I7129,I13341,I14822,g2624,g1569,
    g2373,I15222,g8834,I12271,g3285,g1689,g6966,g8761,I10451,g5216,g5223,
    I13846,g3500,g8172,I14067,I5407,I13731,I5868,g2927,g2677,I14130,I9660,
    g5679,I10172,I11413,I5718,I13704,I10976,I5535,g4584,g6568,g4539,g2881,
    g8746,I14442,g4677,g5831,I10516,g2149,I5894,I6163,I12499,g6597,g7043,g9141,
    I9672,g5576,g6736,I9132,g4284,I6143,I9209,g4349,I12936,I7987,g3528,g5805,
    I10448,g5916,g5022,g4438,g2699,g4019,g6090,g5529,g4362,I11929,g6190,I12989,
    g6932,I6805,g7034,g5749,g5207,I11656,I12340,I14825,g8651,g3523,I14370,
    g7603,I11425,I12722,g6611,g7565,I13865,g2961,I5664,g3643,g2453,I12924,
    g6983,I13583,g7252,I5984,g1564,g642,g7147,I16122,g9353,I10151,g5007,g7347,
    I13457,I15516,g8977,I9558,g4597,g5798,I10433,g7555,g1826,g6663,g7545,
    I10807,I14996,I11371,I8989,g4537,I13779,g3634,I7107,I8193,g3547,g6155,
    I10826,I14844,g8641,I12424,I11392,I11787,g6273,I14394,g7536,I12753,g6445,
    g8866,I15184,g7210,I13144,g3499,I8971,g4464,I12145,g1638,g5796,I7738,g3038,
    g5873,g7164,g5037,I15723,I12199,g6475,g7013,I16049,g5437,g5041,I11827,
    g6231,g7413,I13524,I13743,g7454,g5028,I14420,g7554,I15208,g8810,g2818,
    g1792,g6063,I10678,g6628,g2867,g3754,g2543,g4698,g8198,g8747,g8545,g4025,
    I7792,I14318,g7657,I10236,I12696,g6503,I16148,I14227,g7552,I5689,I7959,
    g2793,g1758,g1589,I14025,g7500,g3578,I11803,g6280,g2470,g9069,I12939,
    I11132,g5917,g7317,I13383,I14058,g7544,g6254,I5428,g6118,g5549,g6167,
    I10862,I11281,g1571,g3983,I11428,g9180,I12487,g7601,g7450,I15607,g8994,
    g9380,g9379,I7389,I9396,g1711,I5555,g2274,g6652,I12161,g4678,g3712,g1952,
    g7855,I12400,I15530,g5786,I10403,I7749,g1827,g2614,g1562,I15484,I14196,
    I11506,I8820,g5364,g5124,g8980,g2325,g2821,I10377,g5188,g1774,I5616,I12708,
    g6482,g7581,I13888,I10739,g5572,g4087,I7882,g4105,I7928,I9076,g5054,g4457,
    I12373,g4801,I9126,I9889,g4819,I14739,g8173,g2348,g3961,g7060,I11890,g6135,
    g1803,g7460,g7172,I6160,g5725,g4465,I11482,g6117,g6598,g3927,I7584,I5609,
    I12244,g6098,I13710,g7340,g2636,I14088,I6767,I11290,g4226,g8386,g8014,
    I5883,g2106,g8975,I15429,g3946,g2306,I6075,I15408,g8896,g8976,g6625,I11867,
    g1662,g2790,g7937,I14285,I7762,g3029,g6607,g6232,I11031,I11778,g6180,g3903,
    I7498,I15690,I12068,I10427,g5210,g7479,I16026,I9850,I10366,g5715,g6253,
    g6938,I14427,g7835,I5466,I13314,I8360,g3513,I9139,g4364,g7190,I13112,g2622,
    g1568,I11945,g5874,I12337,g6724,I5365,I5861,I11356,g7221,g1816,I9639,I8721,
    I13679,I11380,g5822,g5202,g5787,g4007,I7752,g2904,I14403,g7679,g7156,
    I13042,I10582,g6552,I11722,g7356,I13484,g4920,g6606,I11824,g4578,g2917,
    I11090,g2873,I11998,I14657,I7296,I11233,g6147,g2514,g4718,I9018,g8483,
    I8962,I7064,g2458,I11672,g1847,g4803,g9075,g7242,g3743,g2403,g8636,g1685,
    I5528,g2145,g6687,g2345,g2208,g7704,I14001,g4582,g2922,g3916,I7545,g9323,
    g6586,g8790,g2695,g4015,g2637,g1581,I11449,I12918,I10183,g8061,I14330,
    I10292,g8971,I14127,g7594,g7163,I7640,I11897,g6141,I6078,I11961,g7032,
    g2536,I9493,g7354,g8756,g1757,g5309,g7432,I13559,I10786,I12451,g2359,I8907,
    g3560,g2361,g9351,I16103,g2223,I5942,I7844,g3784,I15982,g9236,g5808,I10457,
    g636,I6680,g6645,I11917,I16040,g9285,g4721,I9025,I14103,I11212,g6146,I5852,
    g5759,I10350,g8514,g8040,g3873,g2956,g3095,I6831,g3495,g3653,g2459,I8180,
    I12322,g6751,I14381,g2522,I14181,g7725,g7157,I13045,g2642,g1588,g3936,
    g7357,I13487,g3579,g1929,g3869,I12687,I8853,g4034,I11955,I11401,g6506,
    I11680,g1751,I5847,I12561,g6449,I16183,g9388,g5604,I12295,g6693,g3917,
    I7548,g4670,g1585,g724,g4689,I8966,g6587,I15522,g9018,I15663,g9066,I14190,
    g4279,g6111,g5453,I14448,I11260,g5833,I10522,I7814,g7245,I15959,g4028,
    I7797,g2880,g2234,I7350,g2971,I6864,g2528,I11971,g6179,g4030,g8016,I14311,
    g8757,g5584,g1673,g7712,I15776,I15553,g9009,I13369,I6021,g4564,I8665,
    I11368,g8642,I12364,g6714,g3770,g2551,g5268,I9788,I9014,g5362,I10497,g5233,
    I15536,g9004,g1772,I11467,g4806,g6591,I15702,g9064,I13850,g7328,I12367,
    I5817,g2982,g1848,g3532,I7967,g2787,I14205,g1743,I12430,g2128,g2629,g6020,
    I6127,I10987,g5609,g6702,I5605,I10250,I14076,I8742,g6507,I11683,I8277,
    g1011,I5413,I13228,g6892,I15729,I12253,g6729,I11011,I5751,g5086,I9460,
    g8880,I15218,g3189,I13716,g7475,I13631,I16072,g9303,g3990,g2554,I6376,
    I9681,g4589,I10969,I15672,g7627,I13956,g3888,I15062,g8632,g6905,I12586,
    I13308,g3787,g1842,g8017,g7692,I11880,I15933,g9210,I13758,g5470,g4899,
    I10569,g3956,g5025,I9363,g6515,g6125,I11627,g6630,g4571,g2908,g3675,I7167,
    I12976,g6928,g1573,g1863,I11227,g7021,I13940,I11958,g7039,I9422,I8351,
    I14489,g3811,g2285,g7439,I12643,g6501,I5368,I11386,g5764,I5772,g2490,I6326,
    I6024,I5531,I12669,g6477,g7583,I13894,g7702,I13997,g4196,I10169,I6795,
    g1683,I10503,g5235,g3684,g2180,g3639,g5006,I9333,g3338,I15010,g3963,I7672,
    I15574,g8983,g4538,g2148,I15205,g8809,I6431,g4780,I9089,g1857,I7788,g9050,
    I10177,g5766,I10373,g5087,g1976,I15912,I9095,g4283,I10442,g3808,g7276,
    g5487,I9907,I14315,g7676,g1970,I11793,g6188,I13428,g7167,g3707,g2226,
    I11296,I14819,g8647,I8901,g2698,g4018,I14202,g7708,I8172,g3524,I14257,
    g7716,g4713,g2964,g7495,I16020,g9264,I16161,I7392,g3230,g5755,I15592,g8989,
    I15756,I13761,I14070,g7714,g3957,g6617,I9752,g4705,g4093,I7902,g8512,I8282,
    g3515,I16046,g9288,g1760,g4493,I8543,I11926,I12496,I13822,g3865,g2944,
    I10384,g5193,g6655,g5445,g5059,g3604,I13317,g7211,g5491,g4918,g3498,g7550,
    g7593,g4381,g8649,I14743,g6010,I7302,I11129,g2872,I6590,g1924,I9633,g4685,
    I8952,g4197,I10801,g5463,g6410,I11533,g2734,g4021,I9336,g6968,I14801,g8608,
    g1779,g2057,I12124,I12678,g6516,I12523,I6571,g7120,I9419,I12388,g2457,
    g5578,g5868,I10555,I13388,g2989,g1843,g3539,g3896,I7473,g6143,g5459,I14019,
    g7480,g2393,g5718,I12460,g6674,g7022,I11323,g1977,g7145,g7534,I13299,
    I14695,g7277,I13267,g2834,I6564,I6723,g7220,I14334,g5582,g8902,g6278,g8463,
    g2686,g1667,g7789,I14224,g5261,g2007,I15770,g5793,I10418,I12065,I8202,
    g9332,g6618,g6003,g1665,I10796,I13728,g4562,g6235,I9347,g9199,I16107,I7911,
    g2767,g5218,I8094,g2976,I14457,g8093,g6566,I8808,I13737,g7446,I5359,g8986,
    I13329,I8190,g6134,g5428,g8619,g7547,I13825,I11329,I8264,g5246,I9760,g2625,
    g1570,I8730,g3086,g1852,g2253,g2938,g2347,g3728,g2202,g7433,I13261,g7041,
    g5748,g6555,I11729,g3546,I6946,g1887,I10256,g5401,I12247,I11512,g1732,
    I9675,g4807,I13512,g2969,I5383,I10280,g5488,I14085,g4585,g2925,g6621,
    I11855,g3897,g4041,I11266,g7078,g6683,I13438,I7377,I13831,g7322,I6036,
    I14157,I12277,g6681,g4673,I8928,I10949,I9684,g4813,g7035,g7134,I15803,
    g9148,I7287,g2561,g6094,I10716,I14231,g7566,g4779,I8922,g1565,g649,I8724,
    g5671,I10160,I12782,g6463,I13722,g7442,I16090,g3635,g1949,I13924,I5633,
    g1681,I7781,I6422,g4890,g4075,I12352,g6752,g7280,g2525,I6354,g3801,I7262,
    g7834,I13271,I6419,I8835,g3954,g5826,g6572,g8606,I12170,g4011,I11461,g9076,
    I15622,I5732,g6264,g7310,I13031,g5638,I11407,g2879,I6597,g7025,I11736,
    I11887,I16151,I7344,g2382,g8633,I8799,g3951,g1655,g6050,I12167,g2506,I6437,
    g1784,g6944,I6302,g3091,I13843,g7326,g9267,g3491,g1800,g4080,I7867,g7577,
    g4573,I11764,g6056,g5758,I10347,I13764,I12088,I11365,g2275,g2311,I9539,
    I10896,I13365,g7267,g5466,I10243,g5026,g5624,g7590,I13915,g9184,I15830,
    I13869,g2615,g1563,g4569,g2906,g3920,I12022,g3868,g2174,I11194,I12202,
    I8802,g6224,g2374,I6220,g5448,g5137,g1922,I9162,g4272,g7556,I13161,g7080,
    g5708,g5055,I12313,g6730,I12376,I6733,g5471,g5827,g6585,I12517,I15651,
    g3582,g2284,I5914,g7095,g7064,I12829,g2239,I5978,I7314,g2916,I10180,g9368,
    g1597,g5846,g2380,I6242,I13258,g6907,I12900,g6947,I7870,g2827,g4122,g2184,
    I12466,g5396,g4692,I5636,I12268,I6054,g2020,I5855,I10930,I11043,I6454,
    I12101,I6770,g1590,I11978,g7033,I13861,g8111,I14374,I10387,g4000,I10694,
    I7981,I10965,g6997,g2794,I11069,I15687,I6532,g1694,g9298,g2931,I6669,g3721,
    I7211,g6238,g5027,I13810,g7312,g8174,I15717,g9051,g5467,g4891,g4462,g7194,
    I13118,g7332,I9425,g655,g2905,I6012,g6744,I14064,g8284,I14531,g2628,g3502,
    g7905,I6189,g2630,g5493,g8180,g7719,I14279,g7700,I8739,g4924,I5775,g7966,
    g2100,I7623,I10469,g5222,I11967,I11994,g7471,g7233,g9044,g1942,I6029,g4023,
    I8736,g4008,I10286,I5548,I9669,I15433,g8911,I10552,I6956,g1907,g6901,
    I14039,g7449,g4588,g2929,g5872,g5685,I10186,g5197,I13425,g7166,g4311,g6511,
    I11693,I5398,I15811,g9151,I12454,g6581,g2973,g1854,I5676,g3430,I8910,g4051,
    g3093,g6092,I13918,g9233,I8871,g7150,g6952,I14677,g7791,g7350,I13466,
    I12463,I13444,g7282,g4146,I8011,g7009,I8814,I10937,g5560,I6963,g658,I6109,
    I6791,g1967,g4103,g6721,I8268,I7807,g3910,I7523,I12238,I14178,g2804,I8983,
    g1912,g5631,g7836,I14260,g5723,I9034,g4259,g6772,g3837,g7697,g2351,I6428,
    g3967,I12176,g6510,g8750,I10479,g5227,I12699,g8973,I9369,g7229,g6623,
    I11861,g7993,I14298,I7255,g1955,g5287,I14015,g7440,I9407,I12538,I13656,
    g7228,g3589,I7061,g7699,g5788,g4443,I8449,I13353,g7231,I8477,g9178,I16158,
    g7031,g4116,I12484,I5954,g2884,g2238,I7386,g3048,I6784,I7811,I9582,g4694,
    I8205,g6651,g9182,I5432,g4565,g2901,I14792,g9382,g9217,g8882,g3919,g2372,
    I6214,g7248,I5568,I7341,g2618,g1566,g9355,g2235,I5966,g2343,I10780,I12439,
    g4697,I8986,I11344,g4914,g8178,g2282,I7112,g2546,g1778,g5058,I12385,g4596,
    g3911,g6024,g4013,I12256,g3780,g5129,I12111,g2334,I8273,I12349,g6742,g5722,
    g2548,I7293,I12906,g6918,g8899,g2495,I13023,g7040,g1661,I7329,g2920,I11224,
    g2555,I11028,I11308,g1796,g6711,I15675,I10259,g6523,I11707,I9502,g3972,
    g3994,g4536,I15696,g9208,g9302,g9281,I8862,g6205,I14397,g9074,g2621,g1567,
    I8712,g2712,g1686,I6728,g1959,g5474,g4904,g1646,I8718,I7746,g6634,I11894,
    I13816,g8235,I14492,g2313,I6096,I12120,I5471,g6104,I14964,g8406,I11239,
    I15504,I12138,g4922,g4111,g5439,I13752,g7315,g5844,g2290,g5480,g4913,I6425,
    g1811,g5713,g4581,g3700,I7953,g6754,I12135,g1583,g5569,I8706,I9564,g4703,
    I11669,I13669,g7240,g8792,g5779,g6613,g3950,g4784,g5417,I9053,g5800,I9910,
    g4681,g5688,I10193,I15533,g9002,g2384,I5478,I14747,g8175,I5475,I7716,
    I12457,g4079,I7864,I11525,g6034,g7177,g3562,I7044,I9609,g2264,g6712,g7405,
    I13518,I8919,I6305,g3631,I7098,g7829,g2360,g2933,I6673,g3723,I12609,g6571,
    I13290,I14166,I7198,g2509,g5294,g5000,I5646,g7705,I14807,g8603,g2641,g1587,
    I14974,g8442,I10639,g4501,g2801,g6263,I12684,g3605,g1938,g2996,g1828,I9466,
    g3943,I10353,I15845,I12921,g6993,I13713,g7341,I13250,I8805,g3976,g5468,
    g4195,g1925,g8776,g2724,g1814,g7225,g6936,g7610,I15501,g6014,I10614,I14416,
    g7727,g2379,I13610,g7227,I16145,I12526,g4704,I9001,g6963,g6660,g6946,
    I12649,I13255,g7057,g2878,g2233,I13189,g7002,I7644,g7259,g7124,g6896,
    I12973,g6927,g5608,g4245,I6051,g6903,g2777,g1797,I16009,I10579,g5433,I9774,
    g4250,g2882,I11686,I11939,g6015,I16017,I13460,g4032,I6018,g7275,g7206,
    I13134,I6578,I6868,g6036,I10643,g6913,g1933,I16132,g9356,g5215,I15498,
    g1987,I5842,g4568,g3013,g5665,g5051,I11332,I16043,g3531,g5127,g2674,I11191,
    I11473,g9363,g1776,I7599,I15924,g6767,g4357,g3679,I12286,g5633,g4895,
    I11218,g6161,I5975,g2332,I10430,g5211,I13837,g7324,I7371,g2680,I14430,
    g2353,g4426,g4120,g9183,g6760,g9080,g5696,g1945,I12652,I12265,g1738,g3074,
    I10253,I13305,g3992,I14035,I15199,g5258,g6087,I8793,g3588,I11470,g6095,
    g5240,g5072,g7360,g8799,I14142,g7551,g5472,I9892,g4489,I12490,g7207,I14816,
    g6037,I10646,g3573,I5789,g6102,g8541,g2511,I12478,g1876,g6735,g6064,I11494,
    I13595,g7488,g2092,g5434,g5112,I11037,g7592,g7532,I12131,I13782,g6246,
    g8802,I11419,g1818,g9019,I15481,I7374,g7951,I14288,g3828,I15225,g8689,
    g9072,I10475,I9301,g4295,I12930,I7145,g2501,I5945,I8787,g4475,g3818,g5596,
    g1663,g7870,I14270,g5013,I5709,I14646,I15648,I11215,g2480,g2623,g6725,
    g5706,g5820,I10485,I7359,g2871,g9185,I15833,I7875,g7151,I15657,g9059,g9385,
    I16173,I15068,g8638,I14175,g1877,g5828,g6553,I11725,I15604,I13927,I8745,
    g3929,g2375,g6565,g3220,I15337,I6217,g6012,g1556,g7068,g3779,g4583,g2924,
    g5753,I6039,g6189,g4909,I13749,g7313,g7887,g7122,g3977,I12535,I6048,g5241,
    g5581,I14264,g7698,I9531,g4463,I5911,I6711,g1726,I11440,g8968,I6254,g5060,
    g7352,I11305,g5807,g9331,g6956,g5460,g5597,I11254,I13562,I11981,g6285,
    g4561,g3051,I6333,I9505,g4300,g6664,I15705,g5784,I10397,g4004,g8584,I15918,
    I16033,I10274,I8865,g7496,g4527,g3999,I8856,I7595,g3633,I7104,I6471,I12993,
    g2477,g2643,g6684,g6639,g5668,I11341,g8991,I6509,g4503,I8565,g5840,I7978,
    g2205,g6773,g5190,g4925,g4114,g3732,g2533,g1557,g2634,g3753,I9573,g4701,
    g9045,I15539,g5213,I5401,I14614,g7832,g7266,I13238,g7904,g2104,I5879,I7635,
    I9594,I16023,I7629,g6759,g5524,I13009,g6935,g1948,I15065,g7142,I13012,
    g2926,g9369,I16135,I10565,g5402,g6957,g7255,I8766,g2816,I5380,I14810,g3316,
    I6930,I15571,I11476,g6194,I11596,I7554,g7097,g7497,g5577,g2044,g6604,
    I11818,g5810,I13570,g7198,g6498,g2269,g1773,I8486,I10409,g5204,g4547,g5053,
    I12370,g3987,g3533,g2397,g2862,I15631,g9003,g6682,I9250,g6173,g2039,g9227,
    I15947,g3870,g4838,I6764,g1918,I13241,I9597,g4738,g8754,g6019,I13185,g7020,
    I13092,g7047,I6663,I12514,g6605,g7141,g7129,g8982,g1822,g7329,I13407,g4035,
    I6451,g2946,g2365,I12421,g6486,I14109,g4482,I7964,g3488,g5626,I13921,g3960,
    I9588,I11648,I8105,g3339,I8883,I12098,g9188,I15842,I13157,g9071,g3922,
    g9237,g9216,I12541,g4915,g6156,g6070,g1895,g6897,g1837,I13577,g7186,g6025,
    g7596,g5683,g6755,g4800,g2288,I7118,g2484,g2505,I14091,I6248,g6556,I15669,
    g1768,g7564,I9103,g4374,g7143,g3739,g1698,I6368,I6646,g9171,g3783,g1788,
    g3995,I7728,g3937,g8903,g3079,g5782,I10393,g4002,I10390,g5195,I13906,g7358,
    I13284,g6131,I9443,I7323,g2947,g7149,g2798,g7349,I13463,g7279,g3390,I6949,
    g6766,I10705,I14413,I6856,g4590,g5243,g3501,I13126,I14112,I14267,I15927,
    g2632,g1576,g4297,I8261,g4556,g5084,g5603,g1941,I5812,I6474,g3923,g4317,
    I6443,g7241,I5923,I12760,g6685,g4928,g4119,g6226,g4930,g4121,g8916,g2869,
    g2224,I15610,g8995,g5513,g9048,I5552,g4811,g2389,I7655,I11446,g9060,g2309,
    g9333,g7319,I14904,g8629,g3918,g1958,I6000,I11434,I13472,I13876,g6007,
    I12927,g7014,g9196,g7717,g6059,I12475,g5616,g3568,g1935,g7128,I14712,I6192,
    g6457,I5960,g5200,I13147,g3912,g7686,I7888,g2454,I6294,g2826,g2770,g2210,
    I12250,I10509,g5237,g4557,g2896,I10369,g7599,I15595,g1974,I10933,g8801,
    I10617,g4071,g8752,g6227,I11018,I14851,g8630,I8161,I12965,I8428,I11055,
    I7691,I15160,g8631,I13813,g7314,g8042,g5114,I14623,g6257,g8786,g5120,g6656,
    g9177,g2706,g1821,I8826,g7483,g9194,g3941,I6183,I6608,I10574,g5426,g2371,
    g4200,g1807,I11732,g5617,g8770,g6502,g7710,g5789,I10412,g4009,I16119,g7790,
    g5516,g8990,g6940,I12639,I8308,g7187,I13103,I7311,g5987,g1849,g3778,g7343,
    I5377,g4198,I11491,I9840,g4702,g3735,g6216,g3084,I14305,g6028,I14780,g6646,
    g6671,I14276,g2639,g7046,I12806,g5825,g2216,g2383,g4229,I8140,g5707,g3949,
    I6084,I15693,g9301,I9177,g8029,I7380,g3461,g7345,I13451,g8787,g9282,I7832,
    g2768,I10271,I14160,g3526,I15382,g3998,g5709,g6741,I12117,g8988,I6820,
    g3603,g5478,g7030,I12909,g4921,I7353,g9165,g2957,I8196,g3654,I7931,g2780,
    g1923,g6108,g5435,I11251,g5517,g4258,g5482,g1701,I5545,I12520,g4327,g8684,
    g3583,g4078,g2863,I8775,g8791,I8480,g2498,g6217,g5649,g6758,g6589,I7204,
    I15616,g8997,g2833,I6561,g7251,I13203,g1830,g3952,I7651,g7811,I14238,I8994,
    I10046,g4840,I14046,g7492,g6048,I11991,g2539,I6363,g3561,g9058,I13515,
    g8759,I13882,I12059,g5841,g7271,g1825,g3527,I15385,g6133,g7709,g3647,g5052,
    g2162,I7973,g3071,I6009,I12193,I12629,g3764,g4085,I7878,I7029,g5002,I8847,
    g7595,I13930,I12280,g3503,g3970,I11714,I13441,I12211,I11689,I5670,g1943,
    g1878,I12776,g6739,I13725,g7437,g2728,g2256,g2486,g6018,g7414,I13435,g7170,
    g1934,I11197,I7648,I16154,g3819,g4031,I7804,g7130,g3617,g6093,I11744,g6120,
    g7542,g7330,I11659,I12151,I12319,g5785,g6934,g7355,I8101,g3259,g7783,g3771,
    g1853,I11848,g6159,I9782,g4720,I11398,g5823,I6060,g4286,I10482,g5228,g6700,
    g6244,g6397,I8751,g3892,I9627,g2131,g2006,g2331,g4733,I10545,I13332,g4270,
    g2635,I12659,g8881,g8683,g2105,I7667,g3945,g5452,I12025,g2487,g4358,I9603,
    I14786,g3991,g7090,g4798,I10356,g5711,g8883,g7366,I15519,g5071,g3078,g3340,
    g2474,I10380,g5705,g7056,g6631,g4540,g3590,g5672,I12044,I12085,g7456,g7174,
    I13048,I13767,g3959,g1815,g6101,g7148,I13028,g9161,g7348,g3517,g2283,g3082,
    g9383,I8772,g9220,g9205,g7155,I13481,I12301,g3876,g8131,I14378,g2091,g7273,
    g1960,g5814,g7260,I9576,g3225,I9561,g4695,g8766,g5038,I5395,g3955,I6033,
    g6504,g9358,g7197,g7463,g7239,g5009,g4344,I6286,g7792,g9073,I6299,g8984,
    g4898,g7264,g9127,I15759,I9258,g3516,g5769,I11951,g8755,g5836,g4510,g2840,
    I13234,g7720,I12942,g7367,I12632,I15699,g1676,g2015,g3640,I11431,g3124,
    I12187,I6157,I12403,g6769,I12547,I5989,g7549,I8977,g8999,g1727,g3877,g5212,
    I5692,g8602,g5194,I12226,I13979,g8407,g8013,I7885,g6616,g3657,g4112,g2721,
    g6505,g8868,g7543,g6011,g1746,I14097,g8767,g9043,g3556,I7036,I10343,g5704,
    g3928,g8582,I15738,g6074,g3930,g2502,I6337,g9316,I13541,g7209,g4886,g5716,
    g8015,g7689,I14460,g4879,g5462,g2689,g1670,g6573,I11920,I12980,g6929,I8760,
    g3563,g5205,g6713,g1677,I7658,I12888,g6948,I13828,g7321,I14133,g7574,g691,
    g1866,g2700,I7755,g5475,I7335,I13344,g5537,g4594,g2183,g1855,I12442,I13903,
    g4837,I13173,g7089,g5192,g5085,g3555,I12190,g3966,g2910,g2638,g4065,I7838,
    I14857,g9206,g3677,I14925,g8381,g3948,g4125,g2308,I6081,g7017,g7560,I13755,
    I14009,I7680,g7691,g5642,I13506,g4033,g7087,I14603,g7827,g5520,g1577,g1867,
    I9310,g4268,I7558,I10681,g5686,g5812,I10914,g7158,I6195,g6459,I13490,g6220,
    I11001,I13698,I5386,I15324,I16100,g9338,I12208,g3769,I6952,I14722,I10512,
    g5286,g4714,g1975,I9142,g6977,I7551,g1813,g5538,g6588,g9079,I10842,g2396,
    g3812,I10548,g5260,g6051,g3993,I13770,I9657,g6925,g8793,I6517,g3822,g5610,
    g9005,g5073,g5473,g4081,g6945,I13819,g1872,I9520,g7180,g6103,g7591,g2467,
    g4302,I11395,g5469,g4688,g6696,I9785,g4747,g7420,I11633,I12894,I13701,
    g5206,I13719,g7334,g6508,g6072,g6115,g7678,g1756,I6245,g6274,g8780,I7947,
    g9337,g6009,g5199,g1904,g5747,g5781,g4001,g8018,g8067,I14342,g2263,I13247,
    g6906,I12986,g6931,g8900,g6955,g7054,I11701,g8493,g8041,g5238,g3085,g2781,
    g3485,g1652,g1695,g1637,g4592,g5344,I9819,g6210,g2631,g1586,g4746,I12877,
    g8181,g6596,g2817,g9357,I8998,I12196,g6471,I13140,g6954,I9350,g8421,g5088,
    g4932,g6626,g9082,I9009,g4591,I6959,g3520,g3219,g1687,g2479,g1750,g8076,
    g3958,g7351,g6601,I12866,g8562,g4968,g4576,I15940,I13447,I14709,g6922,
    I5763,I11773,I14680,g6647,g7262,I14199,g3974,g8751,I12223,g2743,g3610,
    g2890,g5245,g5196,g7092,g7701,I15962,g2011,g5806,g3980,g6996,I13776,g4524,
    I12391,g7024,g3540,g9162,g4781,g2074,I5872,I11497,I12885,g7318,g2992,g6165,
    g4577,g2914,g5545,g6686,g3287,I6911,g8772,g1649,I15613,g8996,g4711,g8743,
    g5395,g3898,g4026,g4274,g3510,g6032,g6432,I10454,g7782,g7094,g1823,I13734,
    g4544,I11203,I5542,g7088,g3692,g3694,g8583,g4106,I15507,I7564,g6661,g9320,
    g5481,I12655,g6458,I11377,g5811,g5479,g7160,I13054,I13496,g7179,g4027,
    I5908,g7050,I7632,g6933,g5259,I11870,g5818,I14079,g7579,g6924,g4003,g4676,
    I9496,g3825,g5267,g2161,I8084,g3706,I12502,g4191,g8760,g3008,I8850,g2665,
    g6237,I9845,I10125,g5253,g2327,I6124,g3768,I10783,g5542,g6894,g7269,I13547,
    g4307,g2999,g2346,I6154,g2633,g9244,I10561,g5265,I14687,g5710,I12217,g2157,
    I10295,I15784,g4299,I15628,g9340,g7254,g5592,g7810,g6075,g4016,I12038,
    I6887,g4522,g4115,I7956,g2363,g4552,g1909,g7353,g6603,g7499,g3496,I6974,
    I8877,I7338,g2316,g6283,g5677,I10166,g7335,g3891,I8925,g3913,g3505,g4595,
    g2942,I12666,g6476,g7722,g4341,g4017,g3504,g5198,g4691,g4935,g8993,g1860,
    g8443,g6004,g7826,I11923,g4130,g4542,g3815,g7693,I13088,g9222,g7837,g3497,
    I13885,g9174,I8892,g1879,g4554,g9239,I14668,g7787,g5717,g6949,g7232,I11287,
    g7036,g7561,g5244,I10488,g5230,g9294,g5209,g7476,I8709,g7652,g5264,g3429,
    g4280,I13296,g4512,g2460,I13338,I13287,g2784,g4056,g6959,g5751,g8779,g2937,
    g5752,I13527,g7217,g2668,g8775,g3746,g5083,g7838,g7703,g5566,g8581,g6286,
    g5219,g7077,g5790,g4728,g3953,g5061,g7695,I14294,g7553,g8784,g5461,I13131,
    g7426,g5756,g6035,I11257,g5622,g6276,g5115,g7415,g4057,g3866,g7258,g3716,
    g5514,I6291,g4236,g5191,g8156,g3398,g6110,g7044,g9001,g7983,g7008,g1666,
    g4253,g6643,g5016,g5757,g3644,g8363,I10494,g5232,g7833,g5522,I10466,g2626,
    g3867,g6222,g5654,g5698,g3975,g4586,g6899,g2683,g6930,g6602,g6472,g4570,
    I15645,g4525,g7178,g2782,g5612,I13066,g2627,I14118,I9624,g7443,g6089,g7422,
    g1555,g3680,I13854,g3187,g7625,g6242,g7537,g9252,g4587,g5221,g4275,g8979,
    g3904,g3514,g7037,g6150,g1908,g2276,g9339,g4545,g2616,g5490,g7696,g3359,
    g7436,g2764,g7042,g6262,g4559,g4249,g3757,g6229,g5229,g5217,g3522,g3047,
    g8059,g6281,g3874,g6951,g2521,g2617,g7608,g7412,g7121,g6462,g6215,g8925,
    g7429,g7212,g9144,g9123,g9344,g4123,g8320,I8431,g9259,g8277,I8005,g4351,
    g8299,g6941,g6582,g4410,g8892,g8681,I7994,g5552,g4832,g8945,g6431,g4172,
    I8057,I8058,g7272,g8709,g6176,g6005,g5557,g4343,g8078,g7634,g8340,g6405,
    g4282,g7604,g1714,g5570,g1759,g8690,g4334,g8876,g8769,g6733,g3613,g4804,
    g8915,g8794,g8239,g7419,g7230,g8310,g4494,I8546,I8547,g8824,g8877,g8773,
    g6399,I9330,g9142,g9124,g8928,g5020,g4933,g4320,g8930,I8114,g8064,g4158,
    g4724,g4038,g6440,g4379,g8295,g8237,g6923,g6570,I9222,g8844,I8594,I9166,
    g8089,g7658,g8731,g4271,g5511,g8071,g7540,g8705,g4799,I8033,g8948,g5969,
    g5564,g7602,g6627,g5123,g4132,I8496,g4238,I8157,g8814,g6408,g8150,g4744,
    g3525,g8438,g6972,g5661,g7222,g8836,g4901,g4288,I9261,g6433,g8229,g9349,
    g8822,g6395,g8921,g4417,g5334,g4887,g5548,g4826,g4403,g6266,g8837,g6705,
    g8062,g8620,g8462,g9119,g9049,I8001,g9258,I8401,g4175,g4375,g5313,g4820,
    g6726,g6154,g8842,g7609,g8298,g5094,g9274,g4139,I8000,g4384,g4517,g8854,
    g8941,g4424,g6979,g5095,g5593,g4110,g6112,g5673,g4077,g6001,g5540,g6401,
    g8708,g7575,g5050,g1725,g6727,g8405,g4099,g4304,g8829,g8286,g8798,g8733,
    g8270,g8610,g9345,g4269,I8209,I8524,g8069,g4712,g4276,g6124,g9159,g9138,
    g9359,g8377,g7093,g6673,g4729,g4059,g4961,g9016,g8904,g8287,I8186,g5132,
    I9534,I9535,g8849,I7995,g9251,g4414,I8412,I8413,g3313,g4187,g8291,g3094,
    g1898,g4436,g6142,g4160,g7435,g4378,g4135,g5092,g4182,I8071,I8072,I8240,
    g9272,g8259,g5714,g8088,g8852,g8923,I8461,g6734,g4422,g8701,g9328,g6465,
    g4216,g9130,g9054,g2972,I8046,g8951,g8785,g8314,g4437,g8825,g8650,g1728,
    g8336,g6061,g5257,g8943,g6046,I8115,I8642,g8322,I10597,g8934,g9348,g6145,
    g4054,g3767,g4454,g5077,g4532,I8617,I8618,g6107,g8845,I9202,g8337,g4412,
    g5104,g6757,g9279,g4389,I8612,g6416,I8417,g9118,g9046,g4787,g6047,g8266,
    g6447,g4956,g2979,g1733,g5044,g8081,g8815,g7183,g6132,g4169,g8692,g8726,
    g4138,g4109,g4791,g4707,g4062,g6417,I8090,I8490,g4201,I8108,I8109,g8267,
    g8312,g6629,g6023,g4957,g4049,I8456,I8529,g8293,g8329,g4469,g4889,g4098,
    g6554,g5762,g8828,g8830,g8727,g5436,g6719,I8063,g8703,g8932,g6166,g8624,
    g8953,g8758,g4052,g7687,g4452,g3760,g6456,g6116,g7444,g9158,g9137,g5036,
    g4086,g4179,g4486,I8528,g8716,g7428,g4504,I8568,I8569,g4185,g9275,g4385,
    g8848,g5579,g4090,g4425,g2386,g5442,g4679,g6057,g4131,g8319,I8552,g8258,
    g6971,g6424,g8717,g7597,g7316,g7079,g8274,g4445,I8455,g4091,g4491,g8325,
    g8821,I8052,I8053,g5029,g4369,g8280,g8939,g4407,g4227,g8306,g4793,g3887,
    g8461,g8622,g4246,g3226,g8403,g8841,g5049,I8020,g8695,g8307,g9278,g4388,
    g8359,g9143,g9122,g9343,g7626,g8858,g4430,I8436,I8437,g9334,g8315,g4239,
    g6239,g5314,g5019,g2935,g7683,g4876,g8654,g6420,g4108,g4883,I8040,g4066,
    g8272,g4466,I8491,g8909,g8612,g6204,g4365,g4048,g8935,g5425,g4448,I8460,
    g4072,g8328,g4133,g4333,g8542,g8330,g4396,g9160,g9139,g6040,g5105,g7616,
    g4163,g4067,I8143,g3049,g8090,g6151,g8823,g5045,g5091,g4181,g8456,g9271,
    g4397,g8851,g4421,g8698,g8260,g6172,g9238,g8720,g4101,g8318,g8652,g8843,
    I8593,g8457,g1753,g8686,g4529,g8321,g6908,g4168,g6567,g6265,g4368,g8938,
    g8813,g5030,g4058,g3656,g4743,g3518,g8740,g6965,g6489,g4411,g8687,g6160,
    g1919,g4074,g5108,g6641,g6770,g3678,g5066,g8860,g8341,g8710,g9384,g8645,
    g8691,g5048,g9024,g8884,g8879,g8782,g8154,g8962,g8890,g6249,g1739,g8275,
    g8311,g4400,g3614,g6541,g6144,I8574,g5018,g5067,g5093,g9273,g4147,g4383,
    g4220,g8380,g8832,g4176,g4514,g8853,g7081,g4423,g3188,g5700,g4361,g8931,
    g4127,g4451,g6574,g5984,g7038,g6466,g8628,g8300,g9014,g8906,g7010,g5817,
    g4472,g8440,I8523,g5585,g4741,I8643,g6175,g4332,g5614,g8323,g9335,g4870,
    g4434,I8014,I8015,I8551,g9022,g8887,g4255,g8151,g8648,g6470,g5458,g4686,
    g3509,I8613,g8839,g9037,g8965,g4936,g4117,g8278,g7192,g7026,g8282,g5080,
    g5573,g3011,g8693,g8334,g6044,g6717,g6444,g8621,g4937,g4309,g8313,g4235,
    g4190,g4390,g5126,g9012,g8908,I8288,g4356,g9371,g9352,g6414,g8264,I8041,
    g8933,g7016,g4053,g5588,g3028,g4453,I8495,g6182,g8724,g8379,g7199,g7003,
    g6916,g6022,g5595,g8878,g8777,g6422,g8289,g8835,g8271,g8611,g5043,I8296,
    g6437,g5443,g5116,g8238,g5034,g8332,g4497,g8153,g8744,g7215,g6042,I8029,
    g8804,g6054,g4526,g6615,g2889,g7136,g5117,g8714,g9025,g8889,g4243,g1690,
    g6412,g6688,g6990,g8262,g6171,g5363,g8736,g6429,g6716,g9131,g9055,g8623,
    g7690,g7096,g8722,g7195,g5937,g5562,g5079,g4546,g5141,g8285,g9226,g6109,
    g4224,I8127,g8384,g8339,I8299,g8838,I8019,g8737,g4906,g4789,g2751,g6049,
    g8077,g8643,g6715,g5681,g5032,g5432,g3233,g3358,g9015,g8905,g8742,g8304,
    g8926,g6162,g6268,g7001,g3722,g8273,g6419,g6052,g8269,g4959,I8006,g4435,
    g4690,g4082,g8712,g8543,g8729,g8961,g8885,g9247,g8927,I8045,g5894,g8660,
    g8147,g8946,g7503,g6006,g5575,g3260,g3221,g8513,g6406,g3190,g6105,g4877,
    g8378,g6487,g5750,g8335,g8831,g8288,g8382,g5484,g5096,g8749,g4785,g1678,
    g6045,g5583,g1775,g5712,g8947,g6407,g6578,g6218,g4194,I8089,g8653,g4394,
    g8302,g6600,g8719,g3986,g6415,g5970,g5605,I8028,g8265,g4955,g4254,g4150,
    g2949,g9021,g8886,g8296,g4409,g8725,g6689,g6698,g5547,g1819,g7427,I8589,
    g6428,g6430,g8281,g5078,g6638,g8297,g5082,g8745,g8338,g8963,g8891,g2986,
    g7416,g7140,g8309,I8418,g6448,g6055,g5239,g7654,g4142,g4192,g4392,g6196,
    g4927,g5615,g6396,g8715,g7363,g8833,g6706,g7417,g7144,g8146,g9011,g6418,
    g6994,g3658,g6926,g8268,g5064,g8362,g4958,I8064,g4376,g5070,g1913,g6021,
    g5594,g6421,g8728,g8730,g4225,g8385,g4073,g4796,g8070,g5089,g4473,g4912,
    g4124,g4377,g8331,g9023,g8888,g4287,I8237,g4483,g8087,g8305,g4199,g5438,
    g6041,g5189,g8748,g9327,g4797,g3893,g9146,g9135,g9346,g1834,I8573,g6168,
    g6058,g5561,g7193,g6911,g6743,g8283,g9240,g7682,g8920,g8459,g6411,g8718,
    g7598,g3222,g8261,g6474,g6203,g8637,g6992,g6610,g6694,g4314,I8400,g9147,
    g9136,g5062,g9347,g4228,g8721,g7606,g4408,g9013,g8907,g5298,g4399,g8940,
    I8588,g4230,g6400,g4433,g4427,g5031,g7607,g7325,g8826,g4395,g8741,g5005,
    g6423,g5765,g8609,g7828,g8308,g7615,g3229,g8066,I8034,g4342,g6999,g6633,
    g8711,g5069,g4097,g5343,g8455,g4154,g8827,g8333,g6732,g8846,g6753,g4155,
    g4783,g6043,g4312,g7628,g6434,g8290,g4129,g8256,g4830,g8816,g6914,g6013,
    g5589,g6413,g8700,g7323,g8263,g8950,g4068,I8079,g8723,g8257,g8817,g8301,
    g6060,g4699,g6178,g4398,g5008,g7278,g6995,g6435,g8441,g6699,I8432,g9084,
    g8964,g5830,g5065,g5122,g4319,g4352,g5033,g8458,g4186,g9276,g4386,g5518,
    g8074,g6053,g4083,g8080,g8713,g5142,g6157,g5081,g9120,g9052,I8078,g9277,
    g4387,g8688,g8857,g5783,g7724,g7337,g6121,g8326,g4145,g4391,g5001,g4107,
    g6436,g4159,g8383,g8924,g7611,g4507,g8634,g5483,g4315,g4047,g8361,g4474,
    g6707,g5140,g4166,g8327,g6039,g5068,g6439,g8303,g8696,g8732,g3286,g8944,
    g5699,g7600,g4128,g3081,g1682,g8316,g6970,g5035,g5119,g8697,g8914,g8795,
    g4902,g7175,g6893,g5599,g4745,g4490,g4823,g8820,g4366,g8936,g6771,g8317,
    g5125,g7184,g6138,g4355,g8922,g6738,g8060,g7535,g5106,g6991,g5689,g8460,
    g9038,g8966,g8739,g4055,g4118,g4167,g2783,g4367,g4872,g4549,g8937,g8079,
    g8294,g5046,g8840,g4193,g4393,g6915,g8942,g2912,g5107,g8704,g6002,g5539,
    g6402,g8954,g8763,g6762,g4740,g3258,g5047,g8912,g8796,g6464,g6177,g8929,
    g6728,g7447,g8626,g3984,g5017,g4219,g7182,g6902,g6394,g4962,g6580,g8735,
    g8075,g8949,g7632,g7445,g7653,g8292,g2952,g6438,g4829,g3314,g5090,g8646,
    g6409,g4180,g9270,g4380,g8439,g4420,g4794,g8702,g8919,g8952,g8788,g8276,
    g5063,g4100,g8404,g5118,g8764,g8231,g5057,g3939,g3925,g3915,g3907,I14941,
    g8699,I8225,I15250,I9107,g2214,g8707,g8082,I9047,g6270,I14484,I15055,
    I15051,I15052,I15053,I15054,I15111,g4824,g3315,g8656,I14985,I15019,I15018,
    g3083,g8850,g5040,g3900,g3895,g3890,g4363,g4790,g4786,I15102,I15098,I15099,
    I15100,I15101,g2229,I14771,I15231,I14959,I14960,g8009,I14302,I14951,I14952,
    I15085,g4810,I14759,I15243,I15239,I15240,I15241,I15242,I14758,g4736,I9044,
    g8658,I14990,g4737,g8176,g6452,g2206,g8862,I15169,g8360,g7421,g4318,I15084,
    I15110,g8812,I15254,g2230,I15230,I15265,I15261,I15262,I15263,I15264,I9099,
    I13553,g8819,I14767,g3541,g8811,I15297,I15298,I15041,g5558,I15275,g3602,
    g7062,I14766,I15165,g2014,I15253,I14754,I15175,I15021,I15017,I15020,I15073,
    I15274,g6209,I15292,g8805,g7784,I14219,I14366,I15109,I15283,g6710,I6209,
    g8706,I14980,g8232,I14942,I15040,I15252,I14969,g2213,g3012,g8128,g6910,
    I11603,g6193,g6197,g5556,I15072,I14496,I15152,g8863,I15400,I9029,I15113,
    I15112,g4734,I9038,I14480,I6208,I14468,g8523,g5021,g8694,I15229,I14479,
    I15228,g2995,g8818,I15232,g8680,g8855,I14772,g8847,I14970,g8861,I15031,
    g4735,I9041,g8679,g2262,I15043,I7232,I7233,g4727,g8236,I15284,I15285,
    I14834,I15086,I15082,I15083,g8279,g8613,g8806,g2367,g2352,g2378,g2330,
    I15042,g8859,g7083,I13220,I15030,g6259,g6185,I14933,I15075,I15071,I15074,
    I15276,g8807,g7191,I15272,I15273,g8803,I15251,g3129,g4237,I14932,g6119,
    g8091,g6184,g6174,g6214,g8655,g5546,I14831,I14753,g2368,I5757,I8363,g8230,
    I15290,I15291,I15033,I15029,I15032,g8233,I8224,g2315,g2385,g2294,g2395,
    g2043,I14495,g5555,I14467,I15147,g6153,I15172,g4835,I15044,g8659,I14485,
    I15888,g9192,I15887,I7466,I10092,g4881,I5521,I5519,g4528,I8606,I8607,g5625,
    I7538,I11143,I11142,I7467,g4839,I10906,I12575,I7181,I7179,I11178,I11179,
    I7421,I9548,I9549,I12597,I12598,g4548,I8636,I8637,I15855,I11110,I11108,
    I11177,I6524,I6522,I8510,I8245,I8243,g4313,I11186,I11184,I13685,g7237,
    I6258,I6257,I10889,I10890,I13800,I15819,I15817,I15818,I5600,I5598,I11185,
    I9978,g4880,I9243,g4305,I9241,I6274,I6273,g5284,I10745,I10743,I9746,I9747,
    I9234,g4310,I9233,I6170,I13587,g7234,I6939,g2051,I11117,I11115,g3232,I7531,
    g3938,I7610,I7611,I7505,I7503,I7011,g2333,I7009,I11123,I11122,I11751,
    I11750,g6701,I12032,I12033,I9195,I9196,I13639,g7257,I13638,I10329,I10327,
    I10981,I10982,I6904,g7069,I10328,I10314,I10315,I7480,I7478,I11841,g6158,
    I7569,I7567,I9964,I9963,I7010,g3681,I13786,I13787,I6757,I12051,I6940,I6941,
    I11116,I11615,I11614,I9057,I10991,g5632,I9547,I8255,I8253,g4492,I8537,
    I8538,I7423,I11165,I11163,I6234,I6232,I10744,g5550,I9979,I9980,I10849,
    I10847,I9242,g4476,I8511,I8512,I10790,I10791,I10848,g4871,I7240,I7239,
    g5567,I10361,I10359,I7443,I13600,g7244,I13598,I9691,I10992,I10993,g4231,
    I11137,I11135,I7533,I11873,g6187,I12552,I12550,I9985,g4836,I12870,I12871,
    g9191,I15856,I15857,I6843,I6842,I8119,I8152,I8150,I7460,I7459,I14473,
    I14472,I10789,g5512,I7937,I11136,I7479,I6813,I5599,I10000,I10001,I6740,
    I6739,g4513,I8582,I8583,I11164,I8939,I8938,I13214,I13215,I7156,I8940,
    I11575,I11574,I6997,I6998,I8635,g4831,I11109,I12551,I11102,I11103,I9151,
    g3883,I7453,I7452,I10874,I10875,I7568,I7157,g4869,I8536,I9278,I9276,I7149,
    I7150,I6275,I9235,I10980,I9693,I13640,I10899,I5506,I5507,I11757,g5056,
    g5039,g5023,g6695,I12016,I12017,I7187,I7188,I5520,I10835,I10836,I13397,
    I13395,I6905,I8328,I8326,I6523,I9965,I6750,I13213,g7065,g7082,I10224,
    I10225,I9070,I9071,I10061,g4910,I10060,I7616,g3889,I7437,I7438,I10360,
    I8166,g3231,I8164,I7215,I7216,g4575,I8679,I8680,I15863,I15862,I13396,
    I14246,I14244,I7277,I10071,g4954,I6172,I7617,I12576,I12577,I9153,I13377,
    I13378,I6134,I6133,I12080,I12078,I7892,I7891,I8393,I8392,g1910,I13785,
    I12031,I9476,I9477,I6171,I7140,I7138,I8121,I6202,I6201,I7086,I7087,I12869,
    I6776,I6774,I8605,I7214,I9475,I13003,I13002,I6996,I9692,I6878,I6876,I7180,
    I8659,I8658,I8133,I8134,I12079,I11752,I12596,g5590,I10888,I6103,I6104,
    g4502,I8559,I8560,I10039,I10040,I11149,I8558,I11842,I11843,I7148,I9947,
    I9948,I7436,I12015,I10900,I10901,I9058,I9059,I9946,g4905,I10625,I6135,
    g6559,I6758,I6759,g9202,I15881,I15882,I9182,I9181,I9382,I9381,I10197,
    I10196,I6500,I6499,I10855,I10854,I8151,I13376,I11096,I11094,I10867,I10866,
    I5505,I13802,I10313,g5305,I10819,I10818,I10306,I10307,I11549,g9179,I7085,
    I7485,I6102,I8132,I13686,I13687,I10094,I6203,g4700,I10019,I10017,I10018,
    I11150,I11151,I7270,I7268,I9999,I7609,I9171,g4244,I9169,I10923,I7069,I7068,
    I10300,I10298,I7540,I13004,I10198,I9745,I12853,I12854,I7173,I7174,g9190,
    I15880,I11080,I11078,I6916,I5696,I5695,I7510,I12852,I8503,I8504,I10305,
    I10062,I8678,I7070,I6752,I6917,I5620,I5621,I7241,I5697,I12053,I6233,I10335,
    I10334,I15898,I15899,I14839,I14837,I15897,g9203,I14838,I9069,I10820,g6680,
    g8073,g8092,I11171,I11170,g4893,I10038,I6775,I11079,g5697,I10143,I10142,
    I13599,I10010,I10011,I15850,I15848,I8339,I8338,I9768,I9769,I10093,I11158,
    I11156,I10321,I10322,I11144,I9767,g6722,I10223,I11172,I6539,I6538,I10320,
    I13017,I13016,I11550,I11551,I10953,g5565,I10952,I9170,I7468,I11095,I9826,
    I8660,I10908,I7576,I7574,g4294,I8244,I12052,I9827,I11124,I9152,I13801,
    I8340,I9194,I10834,g5568,I7893,I7186,I11875,I9277,I7444,I7445,I9994,I9992,
    I6751,I7939,I10336,I13018,I7461,I8956,I8955,I6741,I12180,I12181,I13589,
    I13588,g3924,I6066,I6064,I12833,I12834,I11616,I10873,I8957,I7158,I11101,
    I11874,I12832,I10073,I14474,I9828,I8502,g3914,I7532,I12951,I8470,I7512,
    I15889,I9183,I9383,I14245,I7279,I7938,I10144,I8581,I5619,g8644,g4563,
    I10868,I11157,I11576,I10954,I6924,I6923,g6709,I10072,g3894,I10924,I10925,
    I7172,I8165,I9954,I9953,I15864,I10856,I11758,I11759,g5310,g4298,I8254,
    I7575,I9986,I9987,I8120,I6259,g4252,g3906,I7504,I10907,g4911,I7278,I7618,
    I6540,I9993,I7511,I6501,I7139,I7539,I8394,I12952,I12953,g3899,g6163,I12179,
    g4821,I10009,I10627,I8327,I10626,I8472,I15849,I6925,I9955,I10299,I6906,
    g5291,I10080,I10078,I7269,I6877,I7486,I7487,I6844,I7422,g3886,I6814,I10079,
    I6918,g5312,g4359,I7429,I7430,I7454,g4894,g4888,g4884,I7428,g4456,I8471,
    I6065,I6815,g3885,g3310,g8635;

  dff DFF_0(CK,g397,g4635);
  dff DFF_1(CK,g1271,g5176);
  dff DFF_2(CK,g312,g4618);
  dff DFF_3(CK,g273,g4611);
  dff DFF_4(CK,g452,g449);
  dff DFF_5(CK,g948,g8664);
  dff DFF_6(CK,g629,g6827);
  dff DFF_7(CK,g207,g5733);
  dff DFF_8(CK,g1541,g7778);
  dff DFF_9(CK,g1153,g6856);
  dff DFF_10(CK,g940,g5735);
  dff DFF_11(CK,g976,g8864);
  dff DFF_12(CK,g498,g9111);
  dff DFF_13(CK,g314,g4620);
  dff DFF_14(CK,g1092,g7520);
  dff DFF_15(CK,g454,g4639);
  dff DFF_16(CK,g196,g5731);
  dff DFF_17(CK,g535,g3844);
  dff DFF_18(CK,g292,g4613);
  dff DFF_19(CK,g772,g6846);
  dff DFF_20(CK,g1375,g6869);
  dff DFF_21(CK,g689,g6371);
  dff DFF_22(CK,g183,g6309);
  dff DFF_23(CK,g359,g6336);
  dff DFF_24(CK,g1384,g6881);
  dff DFF_25(CK,g1339,g6865);
  dff DFF_26(CK,g20,g6386);
  dff DFF_27(CK,g1424,g3862);
  dff DFF_28(CK,g767,g6841);
  dff DFF_29(CK,g393,g4631);
  dff DFF_30(CK,g1077,g7767);
  dff DFF_31(CK,g1231,g1236);
  dff DFF_32(CK,g294,g4615);
  dff DFF_33(CK,g1477,g9036);
  dff DFF_34(CK,g4,g9372);
  dff DFF_35(CK,g608,g6806);
  dff DFF_36(CK,g1205,g1204);
  dff DFF_37(CK,g465,g6352);
  dff DFF_38(CK,g774,g6848);
  dff DFF_39(CK,g921,g916);
  dff DFF_40(CK,g1304,g1312);
  dff DFF_41(CK,g243,g6318);
  dff DFF_42(CK,g1499,g7772);
  dff DFF_43(CK,g80,g6778);
  dff DFF_44(CK,g1444,g5185);
  dff DFF_45(CK,g1269,g5740);
  dff DFF_46(CK,g600,g6807);
  dff DFF_47(CK,g423,g9105);
  dff DFF_48(CK,g771,g6845);
  dff DFF_49(CK,g803,g7757);
  dff DFF_50(CK,g843,g2647);
  dff DFF_51(CK,g315,g4621);
  dff DFF_52(CK,g455,g4640);
  dff DFF_53(CK,g906,g901);
  dff DFF_54(CK,g622,g6821);
  dff DFF_55(CK,g891,g3855);
  dff DFF_56(CK,g1014,g1012);
  dff DFF_57(CK,g984,g9133);
  dff DFF_58(CK,g117,g5153);
  dff DFF_59(CK,g137,g5150);
  dff DFF_60(CK,g527,g9110);
  dff DFF_61(CK,g1513,g1524);
  dff DFF_62(CK,g278,g6323);
  dff DFF_63(CK,g1378,g6880);
  dff DFF_64(CK,g718,g7753);
  dff DFF_65(CK,g598,g6797);
  dff DFF_66(CK,g1182,g1160);
  dff DFF_67(CK,g1288,g7527);
  dff DFF_68(CK,g1382,g6888);
  dff DFF_69(CK,g179,g5159);
  dff DFF_70(CK,g624,g6831);
  dff DFF_71(CK,g48,g9362);
  dff DFF_72(CK,g362,g9093);
  dff DFF_73(CK,g878,g890);
  dff DFF_74(CK,g270,g9092);
  dff DFF_75(CK,g763,g6836);
  dff DFF_76(CK,g710,g7751);
  dff DFF_77(CK,g730,g7754);
  dff DFF_78(CK,g295,g4616);
  dff DFF_79(CK,g1037,g7519);
  dff DFF_80(CK,g1102,g6855);
  dff DFF_81(CK,g483,g6356);
  dff DFF_82(CK,g775,g7759);
  dff DFF_83(CK,g621,g6819);
  dff DFF_84(CK,g1364,g6878);
  dff DFF_85(CK,g1454,g5187);
  dff DFF_86(CK,g1296,g7304);
  dff DFF_87(CK,g5,g9373);
  dff DFF_88(CK,g1532,g7781);
  dff DFF_89(CK,g587,g3852);
  dff DFF_90(CK,g741,g9386);
  dff DFF_91(CK,g13,g7308);
  dff DFF_92(CK,g606,g6804);
  dff DFF_93(CK,g1012,g6851);
  dff DFF_94(CK,g52,g6781);
  dff DFF_95(CK,g646,g4652);
  dff DFF_96(CK,g1412,g5745);
  dff DFF_97(CK,g327,g6332);
  dff DFF_98(CK,g1189,g6392);
  dff DFF_99(CK,g1389,g4658);
  dff DFF_100(CK,g1029,g2654);
  dff DFF_101(CK,g1371,g6868);
  dff DFF_102(CK,g1429,g2671);
  dff DFF_103(CK,g398,g4636);
  dff DFF_104(CK,g985,g7515);
  dff DFF_105(CK,g354,g4624);
  dff DFF_106(CK,g619,g6817);
  dff DFF_107(CK,g113,g5148);
  dff DFF_108(CK,g133,g5149);
  dff DFF_109(CK,g180,g5158);
  dff DFF_110(CK,g1138,g7524);
  dff DFF_111(CK,g1309,g1308);
  dff DFF_112(CK,g889,g7101);
  dff DFF_113(CK,g390,g6341);
  dff DFF_114(CK,g625,g6823);
  dff DFF_115(CK,g417,g9103);
  dff DFF_116(CK,g681,g7748);
  dff DFF_117(CK,g437,g6348);
  dff DFF_118(CK,g351,g9100);
  dff DFF_119(CK,g1201,g1200);
  dff DFF_120(CK,g109,g6785);
  dff DFF_121(CK,g1049,g8673);
  dff DFF_122(CK,g1098,g6854);
  dff DFF_123(CK,g200,g199);
  dff DFF_124(CK,g240,g6317);
  dff DFF_125(CK,g479,g4649);
  dff DFF_126(CK,g126,g6789);
  dff DFF_127(CK,g596,g6795);
  dff DFF_128(CK,g1268,g5175);
  dff DFF_129(CK,g222,g6313);
  dff DFF_130(CK,g420,g9104);
  dff DFF_131(CK,g3,g9360);
  dff DFF_132(CK,g58,g7734);
  dff DFF_133(CK,g172,g1270);
  dff DFF_134(CK,g387,g6340);
  dff DFF_135(CK,g840,g2648);
  dff DFF_136(CK,g365,g9094);
  dff DFF_137(CK,g1486,g8226);
  dff DFF_138(CK,g1504,g7773);
  dff DFF_139(CK,g1185,g1155);
  dff DFF_140(CK,g1385,g6883);
  dff DFF_141(CK,g583,g3851);
  dff DFF_142(CK,g822,g7512);
  dff DFF_143(CK,g1025,g8871);
  dff DFF_144(CK,g969,g966);
  dff DFF_145(CK,g768,g6842);
  dff DFF_146(CK,g174,g7737);
  dff DFF_147(CK,g685,g7749);
  dff DFF_148(CK,g1087,g6853);
  dff DFF_149(CK,g355,g4625);
  dff DFF_150(CK,g911,g906);
  dff DFF_151(CK,g1226,g6859);
  dff DFF_152(CK,g99,g6783);
  dff DFF_153(CK,g1045,g8224);
  dff DFF_154(CK,g1173,g7526);
  dff DFF_155(CK,g1373,g6871);
  dff DFF_156(CK,g186,g3830);
  dff DFF_157(CK,g760,g6833);
  dff DFF_158(CK,g959,g5169);
  dff DFF_159(CK,g1369,g6875);
  dff DFF_160(CK,g1007,g8867);
  dff DFF_161(CK,g1459,g3863);
  dff DFF_162(CK,g758,g6840);
  dff DFF_163(CK,g480,g6355);
  dff DFF_164(CK,g396,g4634);
  dff DFF_165(CK,g612,g6811);
  dff DFF_166(CK,g38,g5746);
  dff DFF_167(CK,g632,g6830);
  dff DFF_168(CK,g1415,g5180);
  dff DFF_169(CK,g1227,g7108);
  dff DFF_170(CK,g246,g6319);
  dff DFF_171(CK,g449,g3840);
  dff DFF_172(CK,g517,g4651);
  dff DFF_173(CK,g118,g6787);
  dff DFF_174(CK,g138,g6792);
  dff DFF_175(CK,g16,g1404);
  dff DFF_176(CK,g284,g9086);
  dff DFF_177(CK,g142,g6793);
  dff DFF_178(CK,g219,g6312);
  dff DFF_179(CK,g426,g9106);
  dff DFF_180(CK,g1388,g6882);
  dff DFF_181(CK,g806,g7510);
  dff DFF_182(CK,g846,g2646);
  dff DFF_183(CK,g1428,g2672);
  dff DFF_184(CK,g579,g3850);
  dff DFF_185(CK,g1030,g7518);
  dff DFF_186(CK,g614,g6812);
  dff DFF_187(CK,g1430,g4666);
  dff DFF_188(CK,g1247,g6380);
  dff DFF_189(CK,g669,g7745);
  dff DFF_190(CK,g110,g109);
  dff DFF_191(CK,g130,g6790);
  dff DFF_192(CK,g225,g6314);
  dff DFF_193(CK,g281,g9085);
  dff DFF_194(CK,g819,g7761);
  dff DFF_195(CK,g1308,g6385);
  dff DFF_196(CK,g611,g6810);
  dff DFF_197(CK,g631,g6829);
  dff DFF_198(CK,g1217,g6377);
  dff DFF_199(CK,g104,g6784);
  dff DFF_200(CK,g1365,g6867);
  dff DFF_201(CK,g825,g7513);
  dff DFF_202(CK,g1333,g6863);
  dff DFF_203(CK,g474,g4644);
  dff DFF_204(CK,g1396,g4662);
  dff DFF_205(CK,g141,g5151);
  dff DFF_206(CK,g1509,g7774);
  dff DFF_207(CK,g766,g6839);
  dff DFF_208(CK,g1018,g8869);
  dff DFF_209(CK,g588,g9031);
  dff DFF_210(CK,g1467,g8875);
  dff DFF_211(CK,g317,g4623);
  dff DFF_212(CK,g457,g4642);
  dff DFF_213(CK,g486,g6357);
  dff DFF_214(CK,g471,g6354);
  dff DFF_215(CK,g1381,g6887);
  dff DFF_216(CK,g1197,g1196);
  dff DFF_217(CK,g513,g9116);
  dff DFF_218(CK,g1397,g6389);
  dff DFF_219(CK,g533,g530);
  dff DFF_220(CK,g1021,g8870);
  dff DFF_221(CK,g1421,g5179);
  dff DFF_222(CK,g952,g8668);
  dff DFF_223(CK,g1263,g5737);
  dff DFF_224(CK,g580,g6368);
  dff DFF_225(CK,g615,g6813);
  dff DFF_226(CK,g1257,g5738);
  dff DFF_227(CK,g46,g8955);
  dff DFF_228(CK,g402,g6343);
  dff DFF_229(CK,g998,g1005);
  dff DFF_230(CK,g1041,g7765);
  dff DFF_231(CK,g297,g6324);
  dff DFF_232(CK,g954,g8670);
  dff DFF_233(CK,g105,g104);
  dff DFF_234(CK,g145,g5152);
  dff DFF_235(CK,g212,g4601);
  dff DFF_236(CK,g1368,g6874);
  dff DFF_237(CK,g232,g4606);
  dff DFF_238(CK,g990,g7516);
  dff DFF_239(CK,g475,g4645);
  dff DFF_240(CK,g33,g5184);
  dff DFF_241(CK,g951,g8667);
  dff DFF_242(CK,g799,g7756);
  dff DFF_243(CK,g812,g7758);
  dff DFF_244(CK,g567,g6367);
  dff DFF_245(CK,g313,g4619);
  dff DFF_246(CK,g333,g6334);
  dff DFF_247(CK,g168,g7742);
  dff DFF_248(CK,g214,g4603);
  dff DFF_249(CK,g234,g4608);
  dff DFF_250(CK,g652,g646);
  dff DFF_251(CK,g1126,g8674);
  dff DFF_252(CK,g1400,g6390);
  dff DFF_253(CK,g1326,g7306);
  dff DFF_254(CK,g92,g6794);
  dff DFF_255(CK,g309,g6328);
  dff DFF_256(CK,g211,g4600);
  dff DFF_257(CK,g834,g2650);
  dff DFF_258(CK,g231,g4605);
  dff DFF_259(CK,g557,g6366);
  dff DFF_260(CK,g1383,g6889);
  dff DFF_261(CK,g1220,g6378);
  dff DFF_262(CK,g158,g7740);
  dff DFF_263(CK,g627,g6825);
  dff DFF_264(CK,g661,g7743);
  dff DFF_265(CK,g77,g6777);
  dff DFF_266(CK,g831,g2651);
  dff DFF_267(CK,g1327,g7307);
  dff DFF_268(CK,g293,g4614);
  dff DFF_269(CK,g1146,g1612);
  dff DFF_270(CK,g89,g92);
  dff DFF_271(CK,g150,g7738);
  dff DFF_272(CK,g773,g6847);
  dff DFF_273(CK,g859,g8221);
  dff DFF_274(CK,g1240,g1235);
  dff DFF_275(CK,g518,g6361);
  dff DFF_276(CK,g1472,g8960);
  dff DFF_277(CK,g1443,g4667);
  dff DFF_278(CK,g436,g4638);
  dff DFF_279(CK,g405,g6344);
  dff DFF_280(CK,g1034,g8957);
  dff DFF_281(CK,g1147,g1146);
  dff DFF_282(CK,g374,g4627);
  dff DFF_283(CK,g98,g5146);
  dff DFF_284(CK,g563,g9029);
  dff DFF_285(CK,g510,g9115);
  dff DFF_286(CK,g530,g3842);
  dff DFF_287(CK,g215,g4604);
  dff DFF_288(CK,g235,g4609);
  dff DFF_289(CK,g1013,g1014);
  dff DFF_290(CK,g6,g9374);
  dff DFF_291(CK,g55,g7733);
  dff DFF_292(CK,g1317,g5743);
  dff DFF_293(CK,g504,g9113);
  dff DFF_294(CK,g665,g7744);
  dff DFF_295(CK,g544,g6365);
  dff DFF_296(CK,g371,g368);
  dff DFF_297(CK,g62,g7509);
  dff DFF_298(CK,g792,g5162);
  dff DFF_299(CK,g468,g6353);
  dff DFF_300(CK,g815,g7760);
  dff DFF_301(CK,g1460,g4668);
  dff DFF_302(CK,g553,g9028);
  dff DFF_303(CK,g623,g6822);
  dff DFF_304(CK,g501,g9112);
  dff DFF_305(CK,g1190,g8677);
  dff DFF_306(CK,g1390,g4659);
  dff DFF_307(CK,g74,g6776);
  dff DFF_308(CK,g1156,g1081);
  dff DFF_309(CK,g318,g6329);
  dff DFF_310(CK,g458,g4643);
  dff DFF_311(CK,g342,g9097);
  dff DFF_312(CK,g1250,g7111);
  dff DFF_313(CK,g1163,g2655);
  dff DFF_314(CK,g1363,g6877);
  dff DFF_315(CK,g1432,g5183);
  dff DFF_316(CK,g1053,g8873);
  dff DFF_317(CK,g252,g6321);
  dff DFF_318(CK,g330,g6333);
  dff DFF_319(CK,g264,g9090);
  dff DFF_320(CK,g1157,g1156);
  dff DFF_321(CK,g1357,g8675);
  dff DFF_322(CK,g375,g4628);
  dff DFF_323(CK,g68,g6774);
  dff DFF_324(CK,g852,g2644);
  dff DFF_325(CK,g261,g9089);
  dff DFF_326(CK,g516,g4650);
  dff DFF_327(CK,g536,g6363);
  dff DFF_328(CK,g979,g7104);
  dff DFF_329(CK,g778,g7296);
  dff DFF_330(CK,g199,g3832);
  dff DFF_331(CK,g1292,g7302);
  dff DFF_332(CK,g290,g287);
  dff DFF_333(CK,g1084,g7106);
  dff DFF_334(CK,g1439,g5182);
  dff DFF_335(CK,g770,g6844);
  dff DFF_336(CK,g1276,g6384);
  dff DFF_337(CK,g890,g7102);
  dff DFF_338(CK,g1004,g7105);
  dff DFF_339(CK,g1404,g1403);
  dff DFF_340(CK,g93,g5145);
  dff DFF_341(CK,g2,g9361);
  dff DFF_342(CK,g287,g3836);
  dff DFF_343(CK,g560,g6370);
  dff DFF_344(CK,g1224,g6857);
  dff DFF_345(CK,g1320,g7114);
  dff DFF_346(CK,g617,g6815);
  dff DFF_347(CK,g316,g4622);
  dff DFF_348(CK,g336,g9095);
  dff DFF_349(CK,g933,g5166);
  dff DFF_350(CK,g456,g4641);
  dff DFF_351(CK,g345,g9098);
  dff DFF_352(CK,g628,g6826);
  dff DFF_353(CK,g8,g9376);
  dff DFF_354(CK,g887,g7099);
  dff DFF_355(CK,g789,g7297);
  dff DFF_356(CK,g173,g7736);
  dff DFF_357(CK,g550,g9027);
  dff DFF_358(CK,g255,g9087);
  dff DFF_359(CK,g949,g8665);
  dff DFF_360(CK,g1244,g2659);
  dff DFF_361(CK,g620,g6818);
  dff DFF_362(CK,g1435,g5181);
  dff DFF_363(CK,g477,g4647);
  dff DFF_364(CK,g926,g878);
  dff DFF_365(CK,g368,g3838);
  dff DFF_366(CK,g855,g8220);
  dff DFF_367(CK,g1214,g5736);
  dff DFF_368(CK,g1110,g7299);
  dff DFF_369(CK,g1310,g1309);
  dff DFF_370(CK,g296,g4617);
  dff DFF_371(CK,g972,g2653);
  dff DFF_372(CK,g1402,g6391);
  dff DFF_373(CK,g1236,g1240);
  dff DFF_374(CK,g896,g891);
  dff DFF_375(CK,g613,g6820);
  dff DFF_376(CK,g566,g3848);
  dff DFF_377(CK,g1394,g6388);
  dff DFF_378(CK,g1489,g7770);
  dff DFF_379(CK,g883,g921);
  dff DFF_380(CK,g47,g9389);
  dff DFF_381(CK,g971,g5171);
  dff DFF_382(CK,g609,g6808);
  dff DFF_383(CK,g103,g5157);
  dff DFF_384(CK,g1254,g6381);
  dff DFF_385(CK,g556,g3847);
  dff DFF_386(CK,g1409,g5178);
  dff DFF_387(CK,g626,g6824);
  dff DFF_388(CK,g1229,g7110);
  dff DFF_389(CK,g782,g5734);
  dff DFF_390(CK,g237,g6316);
  dff DFF_391(CK,g942,g2652);
  dff DFF_392(CK,g228,g6315);
  dff DFF_393(CK,g706,g7750);
  dff DFF_394(CK,g746,g8956);
  dff DFF_395(CK,g1462,g8678);
  dff DFF_396(CK,g963,g7764);
  dff DFF_397(CK,g129,g5156);
  dff DFF_398(CK,g837,g2649);
  dff DFF_399(CK,g599,g6798);
  dff DFF_400(CK,g1192,g1191);
  dff DFF_401(CK,g828,g7762);
  dff DFF_402(CK,g1392,g6387);
  dff DFF_403(CK,g492,g6359);
  dff DFF_404(CK,g95,g94);
  dff DFF_405(CK,g944,g6372);
  dff DFF_406(CK,g195,g3831);
  dff DFF_407(CK,g1431,g2673);
  dff DFF_408(CK,g1252,g2661);
  dff DFF_409(CK,g356,g6335);
  dff DFF_410(CK,g953,g8669);
  dff DFF_411(CK,g1176,g5172);
  dff DFF_412(CK,g1376,g6890);
  dff DFF_413(CK,g1005,g1004);
  dff DFF_414(CK,g1405,g5744);
  dff DFF_415(CK,g901,g896);
  dff DFF_416(CK,g1270,g1271);
  dff DFF_417(CK,g1225,g6858);
  dff DFF_418(CK,g1073,g9145);
  dff DFF_419(CK,g1324,g7118);
  dff DFF_420(CK,g1069,g9134);
  dff DFF_421(CK,g443,g9101);
  dff DFF_422(CK,g1377,g6891);
  dff DFF_423(CK,g377,g4630);
  dff DFF_424(CK,g618,g6816);
  dff DFF_425(CK,g602,g6800);
  dff DFF_426(CK,g213,g4602);
  dff DFF_427(CK,g233,g4607);
  dff DFF_428(CK,g1199,g6375);
  dff DFF_429(CK,g1399,g3861);
  dff DFF_430(CK,g83,g6779);
  dff DFF_431(CK,g888,g7100);
  dff DFF_432(CK,g573,g9033);
  dff DFF_433(CK,g399,g6342);
  dff DFF_434(CK,g1245,g1244);
  dff DFF_435(CK,g507,g9114);
  dff DFF_436(CK,g547,g9026);
  dff DFF_437(CK,g108,g5147);
  dff DFF_438(CK,g610,g6809);
  dff DFF_439(CK,g630,g6828);
  dff DFF_440(CK,g1207,g5173);
  dff DFF_441(CK,g249,g6320);
  dff DFF_442(CK,g65,g4598);
  dff DFF_443(CK,g916,g911);
  dff DFF_444(CK,g936,g5168);
  dff DFF_445(CK,g478,g4648);
  dff DFF_446(CK,g604,g6802);
  dff DFF_447(CK,g945,g5170);
  dff DFF_448(CK,g1114,g7521);
  dff DFF_449(CK,g100,g99);
  dff DFF_450(CK,g429,g9107);
  dff DFF_451(CK,g809,g7511);
  dff DFF_452(CK,g849,g2645);
  dff DFF_453(CK,g1408,g5177);
  dff DFF_454(CK,g1336,g6864);
  dff DFF_455(CK,g601,g6799);
  dff DFF_456(CK,g122,g6788);
  dff DFF_457(CK,g1065,g9117);
  dff DFF_458(CK,g1122,g8225);
  dff DFF_459(CK,g1228,g7109);
  dff DFF_460(CK,g495,g6360);
  dff DFF_461(CK,g1322,g7116);
  dff DFF_462(CK,g1230,g7300);
  dff DFF_463(CK,g1033,g9034);
  dff DFF_464(CK,g267,g9091);
  dff DFF_465(CK,g1195,g6374);
  dff DFF_466(CK,g1395,g1393);
  dff DFF_467(CK,g373,g4626);
  dff DFF_468(CK,g274,g4612);
  dff DFF_469(CK,g1266,g5739);
  dff DFF_470(CK,g714,g7752);
  dff DFF_471(CK,g734,g7755);
  dff DFF_472(CK,g1142,g8874);
  dff DFF_473(CK,g1342,g7119);
  dff DFF_474(CK,g769,g6843);
  dff DFF_475(CK,g1081,g6852);
  dff DFF_476(CK,g1481,g7769);
  dff DFF_477(CK,g1097,g1185);
  dff DFF_478(CK,g543,g3846);
  dff DFF_479(CK,g1154,g1153);
  dff DFF_480(CK,g1354,g7768);
  dff DFF_481(CK,g489,g6358);
  dff DFF_482(CK,g874,g4654);
  dff DFF_483(CK,g121,g5154);
  dff DFF_484(CK,g591,g9032);
  dff DFF_485(CK,g616,g6814);
  dff DFF_486(CK,g1267,g4656);
  dff DFF_487(CK,g1312,g1311);
  dff DFF_488(CK,g605,g6803);
  dff DFF_489(CK,g182,g5161);
  dff DFF_490(CK,g1401,g1399);
  dff DFF_491(CK,g950,g8666);
  dff DFF_492(CK,g1329,g2663);
  dff DFF_493(CK,g408,g6345);
  dff DFF_494(CK,g871,g5167);
  dff DFF_495(CK,g759,g6832);
  dff DFF_496(CK,g146,g7735);
  dff DFF_497(CK,g202,g5732);
  dff DFF_498(CK,g440,g6349);
  dff DFF_499(CK,g476,g4646);
  dff DFF_500(CK,g184,g6310);
  dff DFF_501(CK,g1149,g7525);
  dff DFF_502(CK,g1398,g1396);
  dff DFF_503(CK,g210,g3834);
  dff DFF_504(CK,g394,g4632);
  dff DFF_505(CK,g86,g6780);
  dff DFF_506(CK,g570,g9030);
  dff DFF_507(CK,g275,g6322);
  dff DFF_508(CK,g303,g6326);
  dff DFF_509(CK,g125,g5155);
  dff DFF_510(CK,g181,g5160);
  dff DFF_511(CK,g1524,g6393);
  dff DFF_512(CK,g595,g576);
  dff DFF_513(CK,g1319,g7113);
  dff DFF_514(CK,g863,g8222);
  dff DFF_515(CK,g1211,g5174);
  dff DFF_516(CK,g966,g8223);
  dff DFF_517(CK,g1186,g1182);
  dff DFF_518(CK,g1386,g6884);
  dff DFF_519(CK,g875,g5165);
  dff DFF_520(CK,g1170,g1173);
  dff DFF_521(CK,g1370,g6876);
  dff DFF_522(CK,g201,g200);
  dff DFF_523(CK,g1325,g7305);
  dff DFF_524(CK,g1280,g7112);
  dff DFF_525(CK,g1106,g7107);
  dff DFF_526(CK,g1061,g9035);
  dff DFF_527(CK,g1387,g6885);
  dff DFF_528(CK,g762,g6835);
  dff DFF_529(CK,g1461,g4669);
  dff DFF_530(CK,g378,g6337);
  dff DFF_531(CK,g1200,g1199);
  dff DFF_532(CK,g1514,g7775);
  dff DFF_533(CK,g1403,g1402);
  dff DFF_534(CK,g1345,g7528);
  dff DFF_535(CK,g1191,g6373);
  dff DFF_536(CK,g1391,g1390);
  dff DFF_537(CK,g185,g4599);
  dff DFF_538(CK,g1307,g3858);
  dff DFF_539(CK,g1159,g1157);
  dff DFF_540(CK,g1223,g6379);
  dff DFF_541(CK,g446,g9102);
  dff DFF_542(CK,g1416,g4665);
  dff DFF_543(CK,g395,g4633);
  dff DFF_544(CK,g764,g6837);
  dff DFF_545(CK,g1251,g6860);
  dff DFF_546(CK,g216,g6311);
  dff DFF_547(CK,g236,g4610);
  dff DFF_548(CK,g205,g3835);
  dff DFF_549(CK,g540,g6364);
  dff DFF_550(CK,g576,g3849);
  dff DFF_551(CK,g1537,g7777);
  dff DFF_552(CK,g727,g8228);
  dff DFF_553(CK,g999,g8865);
  dff DFF_554(CK,g761,g6834);
  dff DFF_555(CK,g1272,g6383);
  dff DFF_556(CK,g1243,g2660);
  dff DFF_557(CK,g1328,g7309);
  dff DFF_558(CK,g1130,g7522);
  dff DFF_559(CK,g1330,g6862);
  dff DFF_560(CK,g114,g6786);
  dff DFF_561(CK,g134,g6791);
  dff DFF_562(CK,g1166,g1167);
  dff DFF_563(CK,g524,g9109);
  dff DFF_564(CK,g1366,g6866);
  dff DFF_565(CK,g348,g9099);
  dff DFF_566(CK,g1148,g1147);
  dff DFF_567(CK,g1348,g7529);
  dff DFF_568(CK,g1155,g1154);
  dff DFF_569(CK,g1260,g6382);
  dff DFF_570(CK,g7,g9375);
  dff DFF_571(CK,g258,g9088);
  dff DFF_572(CK,g521,g6362);
  dff DFF_573(CK,g300,g6325);
  dff DFF_574(CK,g765,g6838);
  dff DFF_575(CK,g1118,g7766);
  dff DFF_576(CK,g1167,g1170);
  dff DFF_577(CK,g1318,g6861);
  dff DFF_578(CK,g1367,g6873);
  dff DFF_579(CK,g677,g7747);
  dff DFF_580(CK,g376,g4629);
  dff DFF_581(CK,g1057,g8959);
  dff DFF_582(CK,g973,g8672);
  dff DFF_583(CK,g1193,g1192);
  dff DFF_584(CK,g1393,g2664);
  dff DFF_585(CK,g1549,g7780);
  dff DFF_586(CK,g1321,g7115);
  dff DFF_587(CK,g1253,g5741);
  dff DFF_588(CK,g1519,g8227);
  dff DFF_589(CK,g584,g6369);
  dff DFF_590(CK,g539,g3845);
  dff DFF_591(CK,g324,g6331);
  dff DFF_592(CK,g432,g9108);
  dff DFF_593(CK,g1158,g1159);
  dff DFF_594(CK,g321,g6330);
  dff DFF_595(CK,g1311,g1310);
  dff DFF_596(CK,g414,g6347);
  dff DFF_597(CK,g1374,g6872);
  dff DFF_598(CK,g94,g6782);
  dff DFF_599(CK,g1284,g7301);
  dff DFF_600(CK,g1545,g7779);
  dff DFF_601(CK,g1380,g6886);
  dff DFF_602(CK,g673,g7746);
  dff DFF_603(CK,g607,g6805);
  dff DFF_604(CK,g306,g6327);
  dff DFF_605(CK,g943,g8671);
  dff DFF_606(CK,g162,g7741);
  dff DFF_607(CK,g411,g6346);
  dff DFF_608(CK,g866,g5163);
  dff DFF_609(CK,g1204,g1203);
  dff DFF_610(CK,g1300,g7303);
  dff DFF_611(CK,g384,g6339);
  dff DFF_612(CK,g339,g9096);
  dff DFF_613(CK,g459,g6350);
  dff DFF_614(CK,g1323,g7117);
  dff DFF_615(CK,g381,g6338);
  dff DFF_616(CK,g1528,g7776);
  dff DFF_617(CK,g1351,g7530);
  dff DFF_618(CK,g597,g6796);
  dff DFF_619(CK,g1372,g6870);
  dff DFF_620(CK,g154,g7739);
  dff DFF_621(CK,g435,g4637);
  dff DFF_622(CK,g970,g963);
  dff DFF_623(CK,g1134,g7523);
  dff DFF_624(CK,g995,g7517);
  dff DFF_625(CK,g190,g201);
  dff DFF_626(CK,g1313,g5742);
  dff DFF_627(CK,g603,g6801);
  dff DFF_628(CK,g1494,g7771);
  dff DFF_629(CK,g462,g6351);
  dff DFF_630(CK,g1160,g1163);
  dff DFF_631(CK,g1360,g8676);
  dff DFF_632(CK,g1450,g5186);
  dff DFF_633(CK,g187,g5730);
  dff DFF_634(CK,g1179,g1186);
  dff DFF_635(CK,g1379,g6879);
  dff DFF_636(CK,g12,g8662);
  dff DFF_637(CK,g71,g6775);
  not NOT_0(g1658,g1313);
  not NOT_1(g1777,g611);
  not NOT_2(I9325,g4242);
  not NOT_3(I7758,g2605);
  not NOT_4(g5652,I10135);
  not NOT_5(I13502,g7135);
  not NOT_6(g6895,I12558);
  not NOT_7(g3880,g2965);
  not NOT_8(g6837,I12382);
  not NOT_9(I15824,g9157);
  not NOT_10(g5843,g5367);
  not NOT_11(I6112,g4);
  not NOT_12(g7189,I13109);
  not NOT_13(g8970,I15414);
  not NOT_14(I6267,g100);
  not NOT_15(g6062,I10675);
  not NOT_16(I16126,g9354);
  not NOT_17(I10519,g5242);
  not NOT_18(I15181,g8734);
  not NOT_19(I11443,g6038);
  not NOT_20(I12436,g6635);
  not NOT_21(I10675,g5662);
  not NOT_22(g2547,I6371);
  not NOT_23(I7365,g3061);
  not NOT_24(I10154,g5109);
  not NOT_25(g1611,g1073);
  not NOT_26(I11278,g5780);
  not NOT_27(g7171,g7071);
  not NOT_28(I14154,g7558);
  not NOT_29(I12274,g6672);
  not NOT_30(g8224,I14451);
  not NOT_31(g5834,I10525);
  not NOT_32(g5971,I10587);
  not NOT_33(g3978,g3160);
  not NOT_34(I6676,g1603);
  not NOT_35(g3612,I7082);
  not NOT_36(I8520,g3652);
  not NOT_37(g2892,g2266);
  not NOT_38(I13469,g7123);
  not NOT_39(I12346,g6737);
  not NOT_40(I9636,g4802);
  not NOT_41(I14637,g8012);
  not NOT_42(g6788,I12235);
  not NOT_43(g1799,I5657);
  not NOT_44(g3935,I7602);
  not NOT_45(I5933,g1158);
  not NOT_46(g9207,g9197);
  not NOT_47(I13039,g6961);
  not NOT_48(I15426,g8895);
  not NOT_49(g5598,g4938);
  not NOT_50(g1674,g1514);
  not NOT_51(g7281,I13277);
  not NOT_52(g3982,g3192);
  not NOT_53(g4666,I8913);
  not NOT_54(I15190,g8685);
  not NOT_55(g2945,g2364);
  not NOT_56(g5121,I9515);
  not NOT_57(g3128,I6839);
  not NOT_58(g3629,g2424);
  not NOT_59(g7297,I13323);
  not NOT_60(g5670,I10157);
  not NOT_61(I11815,g6169);
  not NOT_62(g6842,I12397);
  not NOT_63(g3130,I6849);
  not NOT_64(g9088,I15654);
  not NOT_65(g8789,g8564);
  not NOT_66(g3542,g1777);
  not NOT_67(I12292,g6657);
  not NOT_68(g6298,I11221);
  not NOT_69(g2709,g1747);
  not NOT_70(I11677,g6076);
  not NOT_71(g6392,I11503);
  not NOT_72(g4648,I8859);
  not NOT_73(I8829,g4029);
  not NOT_74(I15546,g9007);
  not NOT_75(g1680,I5515);
  not NOT_76(I15211,g8808);
  not NOT_77(g2340,g1327);
  not NOT_78(I12409,g6398);
  not NOT_79(g4655,I8880);
  not NOT_80(g7745,I14106);
  not NOT_81(g7138,I12996);
  not NOT_82(I6703,g1983);
  not NOT_83(g5938,g5412);
  not NOT_84(g8771,g8564);
  not NOT_85(g2478,g31);
  not NOT_86(g5813,I10472);
  not NOT_87(g7338,I13432);
  not NOT_88(g2907,g2289);
  not NOT_89(g1744,g600);
  not NOT_90(g9215,I15921);
  not NOT_91(g7109,I12915);
  not NOT_92(g6854,I12433);
  not NOT_93(I12635,g6509);
  not NOT_94(g7309,I13359);
  not NOT_95(g1802,g628);
  not NOT_96(I10439,g5214);
  not NOT_97(g2959,g1926);
  not NOT_98(I14728,g8152);
  not NOT_99(I8733,g3996);
  not NOT_100(I14439,g8063);
  not NOT_101(g2517,I6348);
  not NOT_102(g4010,g3097);
  not NOT_103(I7662,g3642);
  not NOT_104(I9446,g3926);
  not NOT_105(I8974,g3871);
  not NOT_106(g5740,I10277);
  not NOT_107(g5519,I9929);
  not NOT_108(g9114,I15732);
  not NOT_109(g1558,I5435);
  not NOT_110(I7290,g2936);
  not NOT_111(g2876,g2231);
  not NOT_112(g9314,I16058);
  not NOT_113(I11884,g6091);
  not NOT_114(I9145,g4264);
  not NOT_115(I6468,g1917);
  not NOT_116(g5606,g4748);
  not NOT_117(I8796,g3934);
  not NOT_118(g7759,I14148);
  not NOT_119(I14349,g7588);
  not NOT_120(I11410,g5845);
  not NOT_121(I12164,g5847);
  not NOT_122(g695,I5392);
  not NOT_123(g6708,g6250);
  not NOT_124(I13410,g7274);
  not NOT_125(I15625,g9000);
  not NOT_126(g6520,I11704);
  not NOT_127(g1901,I5781);
  not NOT_128(g6219,I10998);
  not NOT_129(g6640,I11908);
  not NOT_130(I8980,g4535);
  not NOT_131(g3902,I7495);
  not NOT_132(I12891,g6950);
  not NOT_133(I11479,g6201);
  not NOT_134(I11666,g5772);
  not NOT_135(g5687,I10190);
  not NOT_136(g2915,I6643);
  not NOT_137(I13666,g7238);
  not NOT_138(g6252,g5418);
  not NOT_139(g6812,I12307);
  not NOT_140(g4372,I8357);
  not NOT_141(g7049,I12813);
  not NOT_142(g3512,g1616);
  not NOT_143(I13478,g7126);
  not NOT_144(g5586,g4938);
  not NOT_145(g6958,I12675);
  not NOT_146(I15943,g9214);
  not NOT_147(g4618,I8769);
  not NOT_148(I6716,g1721);
  not NOT_149(g6376,I11455);
  not NOT_150(g4667,I8916);
  not NOT_151(I5981,g459);
  not NOT_152(I8177,g2810);
  not NOT_153(I7847,g3798);
  not NOT_154(I16055,g9291);
  not NOT_155(g9336,I16084);
  not NOT_156(g2310,I6087);
  not NOT_157(g7715,I14022);
  not NOT_158(g1600,g976);
  not NOT_159(g1574,g681);
  not NOT_160(g1864,g162);
  not NOT_161(g4566,g2902);
  not NOT_162(I11556,g6065);
  not NOT_163(g7098,g6525);
  not NOT_164(I5997,g114);
  not NOT_165(g6829,I12358);
  not NOT_166(g7498,I13672);
  not NOT_167(g2663,I6460);
  not NOT_168(I12108,g5939);
  not NOT_169(g6765,I12164);
  not NOT_170(g3529,g2323);
  not NOT_171(g8959,I15391);
  not NOT_172(I6198,g483);
  not NOT_173(g4693,I8974);
  not NOT_174(I13580,g7208);
  not NOT_175(g4134,g3676);
  not NOT_176(g3649,g2424);
  not NOT_177(I14139,g7548);
  not NOT_178(I9416,g4273);
  not NOT_179(I12283,g6692);
  not NOT_180(g8482,g8094);
  not NOT_181(g5525,g4934);
  not NOT_182(g3851,I7356);
  not NOT_183(g5645,g4748);
  not NOT_184(I5353,g3833);
  not NOT_185(g2402,g29);
  not NOT_186(I7950,g2774);
  not NOT_187(g2824,g1688);
  not NOT_188(g1580,g706);
  not NOT_189(g2236,I5969);
  not NOT_190(g7584,I13897);
  not NOT_191(g4555,g2894);
  not NOT_192(g9065,I15589);
  not NOT_193(I9642,g4788);
  not NOT_194(g7539,I13797);
  not NOT_195(I15411,g8897);
  not NOT_196(I15527,g9020);
  not NOT_197(I10415,g5397);
  not NOT_198(I13084,g7071);
  not NOT_199(g9322,g9313);
  not NOT_200(g3964,g3160);
  not NOT_201(g4792,I9111);
  not NOT_202(g9230,I15950);
  not NOT_203(g6225,I11014);
  not NOT_204(I8781,g3932);
  not NOT_205(I8898,g4089);
  not NOT_206(g6073,g5384);
  not NOT_207(g2877,g2232);
  not NOT_208(g6796,I12259);
  not NOT_209(g1736,I5577);
  not NOT_210(I12091,g5988);
  not NOT_211(g4621,I8778);
  not NOT_212(g5607,g4938);
  not NOT_213(g9033,I15513);
  not NOT_214(g7162,I13060);
  not NOT_215(g7268,I13244);
  not NOT_216(g7019,I12771);
  not NOT_217(I11740,g6136);
  not NOT_218(g7362,I13502);
  not NOT_219(g5158,I9600);
  not NOT_220(I13740,g7364);
  not NOT_221(I9654,g4792);
  not NOT_222(I15894,g9195);
  not NOT_223(g6324,I11299);
  not NOT_224(I7723,g3052);
  not NOT_225(g4113,I7950);
  not NOT_226(g6069,I10690);
  not NOT_227(g2556,g1190);
  not NOT_228(g1889,g1018);
  not NOT_229(I7101,g2478);
  not NOT_230(I5901,g52);
  not NOT_231(g2222,I5939);
  not NOT_232(I13676,g7256);
  not NOT_233(g9096,I15678);
  not NOT_234(I8291,g878);
  not NOT_235(I13373,g7270);
  not NOT_236(g2928,g2326);
  not NOT_237(g4202,g2810);
  not NOT_238(g8663,I14783);
  not NOT_239(I7605,g2752);
  not NOT_240(I15714,g9077);
  not NOT_241(g5587,g4938);
  not NOT_242(g2930,g2328);
  not NOT_243(I15315,g8738);
  not NOT_244(I11800,g6164);
  not NOT_245(g1871,I5754);
  not NOT_246(g4908,g4088);
  not NOT_247(g6377,I11458);
  not NOT_248(g6206,g5639);
  not NOT_249(g5311,g4938);
  not NOT_250(g2899,g2272);
  not NOT_251(g9195,I15871);
  not NOT_252(g4094,I7905);
  not NOT_253(I11936,g5918);
  not NOT_254(g3872,g2954);
  not NOT_255(I15202,g8797);
  not NOT_256(g3652,I7132);
  not NOT_257(g4567,g2903);
  not NOT_258(g7728,I14055);
  not NOT_259(g7486,I13646);
  not NOT_260(g3843,I7332);
  not NOT_261(g3989,g3131);
  not NOT_262(I6186,g138);
  not NOT_263(g7730,I14061);
  not NOT_264(I9612,g4776);
  not NOT_265(I10608,g5701);
  not NOT_266(g5174,I9648);
  not NOT_267(g8762,g8585);
  not NOT_268(g7504,I13692);
  not NOT_269(I15978,g9235);
  not NOT_270(I14115,g7563);
  not NOT_271(g7185,I13099);
  not NOT_272(g4776,I9081);
  not NOT_273(I7041,g2401);
  not NOT_274(g6849,I12418);
  not NOT_275(I9935,g4812);
  not NOT_276(g4593,g2939);
  not NOT_277(I11964,g5971);
  not NOT_278(g3549,g2404);
  not NOT_279(g3834,I7305);
  not NOT_280(g3971,I7688);
  not NOT_281(g7070,g6562);
  not NOT_282(g2295,g995);
  not NOT_283(I14052,g7494);
  not NOT_284(g2237,I5972);
  not NOT_285(g7470,g7253);
  not NOT_286(I15741,g9083);
  not NOT_287(g8657,I14763);
  not NOT_288(g6781,I12214);
  not NOT_289(g7425,I13550);
  not NOT_290(g5180,I9666);
  not NOT_291(g2844,I6574);
  not NOT_292(I8215,g3577);
  not NOT_293(g6898,I12567);
  not NOT_294(g1838,g1450);
  not NOT_295(g5591,g4841);
  not NOT_296(g6900,I12571);
  not NOT_297(g8222,I14445);
  not NOT_298(I8886,g4308);
  not NOT_299(g5832,I10519);
  not NOT_300(I14813,g8640);
  not NOT_301(g1795,I5649);
  not NOT_302(g6797,I12262);
  not NOT_303(g1737,g597);
  not NOT_304(g2394,I6270);
  not NOT_305(g9248,I15978);
  not NOT_306(g1809,g759);
  not NOT_307(I10973,g5726);
  not NOT_308(I14798,g8605);
  not NOT_309(g6245,g5690);
  not NOT_310(g4360,I8333);
  not NOT_311(I7368,g3018);
  not NOT_312(g9255,I15985);
  not NOT_313(g9081,I15635);
  not NOT_314(I12948,g6919);
  not NOT_315(I13909,g7339);
  not NOT_316(I15735,g9078);
  not NOT_317(g4521,g2866);
  not NOT_318(I14184,g7726);
  not NOT_319(g1672,g1499);
  not NOT_320(I14674,g7788);
  not NOT_321(g8464,g8039);
  not NOT_322(g6291,I11200);
  not NOT_323(I12702,g6497);
  not NOT_324(g2557,g940);
  not NOT_325(g4050,g3080);
  not NOT_326(g4641,I8838);
  not NOT_327(I11908,g5918);
  not NOT_328(I12757,g6577);
  not NOT_329(g9097,I15681);
  not NOT_330(g2966,g1856);
  not NOT_331(g5794,I10421);
  not NOT_332(I5889,g83);
  not NOT_333(g1643,g1211);
  not NOT_334(I11569,g6279);
  not NOT_335(g7131,g6976);
  not NOT_336(g6344,I11359);
  not NOT_337(g2471,I6309);
  not NOT_338(g7006,I12748);
  not NOT_339(g7331,I13413);
  not NOT_340(I15196,g8778);
  not NOT_341(I6636,g1704);
  not NOT_342(I14732,g8155);
  not NOT_343(g2242,g985);
  not NOT_344(g6207,I10962);
  not NOT_345(g3909,I7520);
  not NOT_346(I11747,g6123);
  not NOT_347(I12564,g6720);
  not NOT_348(g8563,I14662);
  not NOT_349(g2948,g2366);
  not NOT_350(I11242,g6183);
  not NOT_351(g7766,I14169);
  not NOT_352(g6819,I12328);
  not NOT_353(g7105,I12903);
  not NOT_354(g3519,g2185);
  not NOT_355(I10761,g5302);
  not NOT_356(g7305,I13347);
  not NOT_357(I7856,g3805);
  not NOT_358(I7734,g2595);
  not NOT_359(g2955,I6703);
  not NOT_360(g7487,I13649);
  not NOT_361(g5628,g4748);
  not NOT_362(g1742,g1486);
  not NOT_363(g6088,I10708);
  not NOT_364(g6852,I12427);
  not NOT_365(g5515,g4923);
  not NOT_366(I12397,g6764);
  not NOT_367(g6488,I11652);
  not NOT_368(g4658,I8889);
  not NOT_369(g7748,I14115);
  not NOT_370(g4777,I9084);
  not NOT_371(I10400,g5201);
  not NOT_372(g5100,I9484);
  not NOT_373(I9512,g3985);
  not NOT_374(I13807,g7320);
  not NOT_375(I11974,g5956);
  not NOT_376(I12062,g5988);
  not NOT_377(I14400,g7677);
  not NOT_378(g2350,I6166);
  not NOT_379(g9112,I15726);
  not NOT_380(g7755,I14136);
  not NOT_381(g9218,I15930);
  not NOT_382(g1926,g874);
  not NOT_383(I9823,g5138);
  not NOT_384(g9312,I16052);
  not NOT_385(g2038,g809);
  not NOT_386(g4882,g4069);
  not NOT_387(I14214,g7576);
  not NOT_388(I12933,g7018);
  not NOT_389(I9366,g4350);
  not NOT_390(g7226,g6937);
  not NOT_391(I11230,g6140);
  not NOT_392(I11293,g5824);
  not NOT_393(I10207,g5075);
  not NOT_394(I13293,g7159);
  not NOT_395(I12508,g6593);
  not NOT_396(I11638,g5847);
  not NOT_397(g6886,I12529);
  not NOT_398(I6446,g1812);
  not NOT_399(g4611,I8748);
  not NOT_400(g291,I5356);
  not NOT_401(I14005,g7434);
  not NOT_402(g7045,g6490);
  not NOT_403(I11416,g5829);
  not NOT_404(I10538,g5255);
  not NOT_405(I6003,g228);
  not NOT_406(I9148,g4354);
  not NOT_407(I13416,g7165);
  not NOT_408(I5795,g1236);
  not NOT_409(g9129,I15765);
  not NOT_410(g2769,g2424);
  not NOT_411(g7173,g6980);
  not NOT_412(g9329,g9317);
  not NOT_413(g6314,I11269);
  not NOT_414(g7091,g6525);
  not NOT_415(g7491,I13653);
  not NOT_416(g6870,I12481);
  not NOT_417(g3860,I7383);
  not NOT_418(g2918,g2310);
  not NOT_419(g3341,I6936);
  not NOT_420(g1983,I5839);
  not NOT_421(g6825,I12346);
  not NOT_422(g6650,g6213);
  not NOT_423(g7169,I13075);
  not NOT_424(g7283,I13281);
  not NOT_425(g1572,g673);
  not NOT_426(g8955,I15379);
  not NOT_427(I6695,g2246);
  not NOT_428(g4541,g2883);
  not NOT_429(g7059,g6538);
  not NOT_430(g7920,I14282);
  not NOT_431(g7578,I13879);
  not NOT_432(g6008,g5367);
  not NOT_433(I11835,g6181);
  not NOT_434(g3691,I7195);
  not NOT_435(I11014,g5621);
  not NOT_436(g7459,I13617);
  not NOT_437(g9221,I15937);
  not NOT_438(I12205,g6488);
  not NOT_439(I9463,g3942);
  not NOT_440(g7718,I14031);
  not NOT_441(g7767,I14172);
  not NOT_442(g4153,I8024);
  not NOT_443(g4680,I8945);
  not NOT_444(I7688,g3650);
  not NOT_445(g6136,I10773);
  not NOT_446(g4353,g3665);
  not NOT_447(I11586,g6256);
  not NOT_448(I12912,g7006);
  not NOT_449(g6336,I11335);
  not NOT_450(I14100,g7580);
  not NOT_451(I6223,g330);
  not NOT_452(g8038,g7694);
  not NOT_453(g6768,I12173);
  not NOT_454(I8913,g4306);
  not NOT_455(g7582,I13891);
  not NOT_456(g6594,I11796);
  not NOT_457(g1961,g1345);
  not NOT_458(g3879,g2963);
  not NOT_459(g4802,I9129);
  not NOT_460(g7261,I13225);
  not NOT_461(I14683,g7825);
  not NOT_462(g3962,g3131);
  not NOT_463(g5151,I9579);
  not NOT_464(g7793,I14234);
  not NOT_465(g3158,I6853);
  not NOT_466(g3659,g2293);
  not NOT_467(g6806,I12289);
  not NOT_468(g5648,g4748);
  not NOT_469(I6416,g1794);
  not NOT_470(g3506,g1781);
  not NOT_471(g7015,I12763);
  not NOT_472(I12592,g1008);
  not NOT_473(g4558,g2897);
  not NOT_474(g9068,I15598);
  not NOT_475(I7126,g2494);
  not NOT_476(I5926,g297);
  not NOT_477(I7400,g3075);
  not NOT_478(I8859,g3968);
  not NOT_479(I7326,g2940);
  not NOT_480(I6115,g134);
  not NOT_481(I6251,g489);
  not NOT_482(g2921,g2312);
  not NOT_483(g6065,I10684);
  not NOT_484(g6887,I12532);
  not NOT_485(g6122,I10752);
  not NOT_486(I10882,g5600);
  not NOT_487(g6228,I11021);
  not NOT_488(I5754,g966);
  not NOT_489(g3587,g1964);
  not NOT_490(g6322,I11293);
  not NOT_491(I11275,g5768);
  not NOT_492(I9457,g3940);
  not NOT_493(g8918,I15340);
  not NOT_494(I16180,g9387);
  not NOT_495(g6230,I11025);
  not NOT_496(g7246,I13196);
  not NOT_497(g8967,I15405);
  not NOT_498(I13746,g7311);
  not NOT_499(I13493,g7132);
  not NOT_500(I9393,g4266);
  not NOT_501(g4511,g2841);
  not NOT_502(I15660,g9062);
  not NOT_503(g2895,g2268);
  not NOT_504(g6033,g5384);
  not NOT_505(g2837,g1780);
  not NOT_506(g7721,g7344);
  not NOT_507(g5839,I10532);
  not NOT_508(I9834,g4782);
  not NOT_509(g4092,I7899);
  not NOT_510(I13035,g6964);
  not NOT_511(g3985,I7712);
  not NOT_512(I12731,g6579);
  not NOT_513(I11806,g6275);
  not NOT_514(g4600,I8715);
  not NOT_515(I7383,g3465);
  not NOT_516(g4574,g3466);
  not NOT_517(g6096,g5317);
  not NOT_518(g6496,I11662);
  not NOT_519(g1679,I5512);
  not NOT_520(I8097,g3237);
  not NOT_521(g5172,I9642);
  not NOT_522(g5278,I9794);
  not NOT_523(g6845,I12406);
  not NOT_524(g7502,I13682);
  not NOT_525(I15550,g9008);
  not NOT_526(g9198,g9187);
  not NOT_527(g3545,g2344);
  not NOT_528(I8354,g1163);
  not NOT_529(g738,I5404);
  not NOT_530(g6195,I10940);
  not NOT_531(g5618,g5015);
  not NOT_532(g6137,I10776);
  not NOT_533(g6891,I12544);
  not NOT_534(g5143,I9555);
  not NOT_535(g1831,g689);
  not NOT_536(g6337,I11338);
  not NOT_537(g3591,g1789);
  not NOT_538(g3832,I7299);
  not NOT_539(g4580,g2919);
  not NOT_540(g9241,I15971);
  not NOT_541(I7588,g2584);
  not NOT_542(g3853,I7362);
  not NOT_543(I14725,g8145);
  not NOT_544(g7188,I13106);
  not NOT_545(g5988,I10592);
  not NOT_546(g2842,g2209);
  not NOT_547(I9938,g4878);
  not NOT_548(I10758,g5662);
  not NOT_549(g1805,I5667);
  not NOT_550(g6807,I12292);
  not NOT_551(g1916,g775);
  not NOT_552(g5693,I10204);
  not NOT_553(g7216,I13152);
  not NOT_554(g1749,g371);
  not NOT_555(g2298,I6072);
  not NOT_556(I14082,g7539);
  not NOT_557(g6859,I12448);
  not NOT_558(g2392,g11);
  not NOT_559(I13193,g7007);
  not NOT_560(g2485,g62);
  not NOT_561(I11362,g5821);
  not NOT_562(g7028,g6525);
  not NOT_563(I13362,g7265);
  not NOT_564(g3931,I7592);
  not NOT_565(I8218,g3002);
  not NOT_566(I15773,g9126);
  not NOT_567(I6629,g2052);
  not NOT_568(g4623,I8784);
  not NOT_569(g7247,I13199);
  not NOT_570(g1798,I5654);
  not NOT_571(I6130,g560);
  not NOT_572(g4076,I7859);
  not NOT_573(g9319,g9309);
  not NOT_574(I10940,g5489);
  not NOT_575(g2941,g2349);
  not NOT_576(I9606,g4687);
  not NOT_577(g6342,I11353);
  not NOT_578(g3905,g3192);
  not NOT_579(I13475,g7125);
  not NOT_580(g5621,g4748);
  not NOT_581(I14848,g8625);
  not NOT_582(g6255,I11066);
  not NOT_583(g6815,I12316);
  not NOT_584(I10804,g5526);
  not NOT_585(I6800,g2016);
  not NOT_586(I9687,g4822);
  not NOT_587(g3630,I7095);
  not NOT_588(g6481,I11641);
  not NOT_589(I14804,g8563);
  not NOT_590(g7741,I14094);
  not NOT_591(g4651,I8868);
  not NOT_592(g5113,I9499);
  not NOT_593(g6692,I12008);
  not NOT_594(g6097,g5345);
  not NOT_595(I11437,g5801);
  not NOT_596(I15839,g9168);
  not NOT_597(g2520,g41);
  not NOT_598(I15930,g9209);
  not NOT_599(g2640,g1584);
  not NOT_600(g9211,I15909);
  not NOT_601(g6354,I11389);
  not NOT_602(g4285,I8233);
  not NOT_603(I8727,g3944);
  not NOT_604(g9186,I15836);
  not NOT_605(I5679,g911);
  not NOT_606(g4500,g2832);
  not NOT_607(g9386,I16176);
  not NOT_608(g6960,I12681);
  not NOT_609(I15965,g9219);
  not NOT_610(I7944,g3774);
  not NOT_611(g1579,g703);
  not NOT_612(g1869,g74);
  not NOT_613(g7108,I12912);
  not NOT_614(I10135,g4960);
  not NOT_615(g7308,I13356);
  not NOT_616(I11347,g5761);
  not NOT_617(g2958,g2377);
  not NOT_618(I13347,g7224);
  not NOT_619(g9026,I15492);
  not NOT_620(I5831,g1194);
  not NOT_621(g2376,I6226);
  not NOT_622(g5494,I9918);
  not NOT_623(g3750,g2177);
  not NOT_624(I9570,g4696);
  not NOT_625(I10406,g5203);
  not NOT_626(I9341,g4251);
  not NOT_627(I10962,g5719);
  not NOT_628(g1752,g603);
  not NOT_629(I14406,g7681);
  not NOT_630(g3973,g3097);
  not NOT_631(I9525,g4413);
  not NOT_632(I11781,g6284);
  not NOT_633(I12768,g6718);
  not NOT_634(I15619,g8998);
  not NOT_635(g9370,I16138);
  not NOT_636(g1917,I5795);
  not NOT_637(I9645,g4900);
  not NOT_638(I15557,g9010);
  not NOT_639(g2829,g1785);
  not NOT_640(g9125,I15753);
  not NOT_641(g4024,g3160);
  not NOT_642(I11236,g6148);
  not NOT_643(g2286,I6042);
  not NOT_644(g6783,I12220);
  not NOT_645(g7758,I14145);
  not NOT_646(g7066,I12839);
  not NOT_647(I10500,g5234);
  not NOT_648(I16168,g9381);
  not NOT_649(g7589,I13912);
  not NOT_650(I6090,g390);
  not NOT_651(g2911,g2292);
  not NOT_652(g4795,I9116);
  not NOT_653(I8932,g4096);
  not NOT_654(I5422,g1234);
  not NOT_655(g7466,I13622);
  not NOT_656(g4809,I9148);
  not NOT_657(g6267,I11086);
  not NOT_658(g6312,I11263);
  not NOT_659(g3969,g3192);
  not NOT_660(I6166,g480);
  not NOT_661(I14049,g7493);
  not NOT_662(g9280,I16006);
  not NOT_663(I11821,g6170);
  not NOT_664(I12881,g6478);
  not NOT_665(g1786,g623);
  not NOT_666(g7365,I13509);
  not NOT_667(g7048,I12810);
  not NOT_668(I7347,g2985);
  not NOT_669(g9083,I15641);
  not NOT_670(g2270,I6015);
  not NOT_671(g4477,I8517);
  not NOT_672(g7448,I13605);
  not NOT_673(I13063,g6973);
  not NOT_674(g7711,I14012);
  not NOT_675(g4523,g2868);
  not NOT_676(g6676,I11984);
  not NOT_677(I11790,g6282);
  not NOT_678(g6293,I11206);
  not NOT_679(I13264,g7061);
  not NOT_680(I6148,g5);
  not NOT_681(g7055,g6517);
  not NOT_682(g8219,I14436);
  not NOT_683(g4643,I8844);
  not NOT_684(g3666,g2134);
  not NOT_685(I9158,g4256);
  not NOT_686(I13137,g7027);
  not NOT_687(I6348,g1354);
  not NOT_688(g2225,I5948);
  not NOT_689(g6129,I10758);
  not NOT_690(g8640,I14728);
  not NOT_691(g7455,I13613);
  not NOT_692(g6329,I11314);
  not NOT_693(g6761,I12154);
  not NOT_694(g2073,g1254);
  not NOT_695(g5160,I9606);
  not NOT_696(g7133,I12983);
  not NOT_697(I7697,g3052);
  not NOT_698(g9106,I15708);
  not NOT_699(g7333,I13419);
  not NOT_700(I13873,g7342);
  not NOT_701(g9306,I16036);
  not NOT_702(g6828,I12355);
  not NOT_703(g1770,g606);
  not NOT_704(g7774,I14193);
  not NOT_705(g5521,g4929);
  not NOT_706(g8958,I15388);
  not NOT_707(g6830,I12361);
  not NOT_708(g4634,I8817);
  not NOT_709(g3648,g2424);
  not NOT_710(g3875,g2958);
  not NOT_711(g2324,I6115);
  not NOT_712(g3530,g2185);
  not NOT_713(I9111,g4232);
  not NOT_714(g7196,I13122);
  not NOT_715(g4742,I9064);
  not NOT_716(g9061,I15577);
  not NOT_717(I15601,g8992);
  not NOT_718(g9187,I15839);
  not NOT_719(g4104,I7925);
  not NOT_720(I10605,g5440);
  not NOT_721(I11422,g5842);
  not NOT_722(g6592,I11790);
  not NOT_723(g3655,g1844);
  not NOT_724(I15187,g8682);
  not NOT_725(I14273,g7631);
  not NOT_726(I11209,g6139);
  not NOT_727(I13422,g7131);
  not NOT_728(I14106,g7586);
  not NOT_729(I13209,g6912);
  not NOT_730(g2540,g1339);
  not NOT_731(I9615,g4739);
  not NOT_732(g6221,I11004);
  not NOT_733(I12003,g6202);
  not NOT_734(g8765,g8524);
  not NOT_735(g7538,I13794);
  not NOT_736(I13834,g7466);
  not NOT_737(I6463,g1769);
  not NOT_738(I10463,g5220);
  not NOT_739(I16084,g9324);
  not NOT_740(g2177,g1322);
  not NOT_741(g7780,I14211);
  not NOT_742(g9027,I15495);
  not NOT_743(g5724,g4969);
  not NOT_744(g2377,I6229);
  not NOT_745(I14463,g8072);
  not NOT_746(I12779,g6740);
  not NOT_747(g5179,I9663);
  not NOT_748(g6703,I12041);
  not NOT_749(g7509,I13707);
  not NOT_750(g4926,g4202);
  not NOT_751(I15937,g9212);
  not NOT_752(g9200,g9189);
  not NOT_753(I11021,g5627);
  not NOT_754(I14234,g7614);
  not NOT_755(g3884,I7417);
  not NOT_756(g3839,I7320);
  not NOT_757(g2287,I6045);
  not NOT_758(g7018,I12768);
  not NOT_759(g4273,I8215);
  not NOT_760(g7067,g6658);
  not NOT_761(g8974,I15426);
  not NOT_762(I7317,g2893);
  not NOT_763(g5658,g4748);
  not NOT_764(I15791,g9140);
  not NOT_765(g7418,I13533);
  not NOT_766(g6624,I11864);
  not NOT_767(g7467,g7236);
  not NOT_768(g6953,g6745);
  not NOT_769(I6118,g243);
  not NOT_770(I14795,g8604);
  not NOT_771(g8225,I14454);
  not NOT_772(g5835,I10528);
  not NOT_773(g7290,I13302);
  not NOT_774(g4613,I8754);
  not NOT_775(g6068,I10687);
  not NOT_776(g1888,g781);
  not NOT_777(I6872,g2185);
  not NOT_778(g9145,I15791);
  not NOT_779(g4044,g2595);
  not NOT_780(g6468,I11622);
  not NOT_781(I12945,g7066);
  not NOT_782(I9591,g4710);
  not NOT_783(g4444,I8452);
  not NOT_784(g1787,g625);
  not NOT_785(I6652,g2016);
  not NOT_786(I11607,g5767);
  not NOT_787(I6057,g518);
  not NOT_788(I12826,g6441);
  not NOT_789(I12999,g7029);
  not NOT_790(I11320,g5797);
  not NOT_791(I15666,g9070);
  not NOT_792(I13320,g7139);
  not NOT_793(I6457,g1886);
  not NOT_794(g7493,I13659);
  not NOT_795(g1675,g1519);
  not NOT_796(g6677,I11987);
  not NOT_797(g7256,g7058);
  not NOT_798(I13274,g6917);
  not NOT_799(I7775,g3705);
  not NOT_800(g5611,g4969);
  not NOT_801(g8324,I14573);
  not NOT_802(g4572,g2909);
  not NOT_803(I7922,g3462);
  not NOT_804(g2898,g2271);
  not NOT_805(I15478,g8910);
  not NOT_806(g2900,g2273);
  not NOT_807(g6866,I12469);
  not NOT_808(I12672,g6473);
  not NOT_809(I7581,g3612);
  not NOT_810(I13122,g7070);
  not NOT_811(g9107,I15711);
  not NOT_812(g4543,g2885);
  not NOT_813(I10421,g5208);
  not NOT_814(I11464,g6088);
  not NOT_815(g5799,I10436);
  not NOT_816(I13565,g7181);
  not NOT_817(I9794,g4778);
  not NOT_818(I6834,g287);
  not NOT_819(g9307,g9300);
  not NOT_820(g2510,g58);
  not NOT_821(g639,I5374);
  not NOT_822(g2245,g999);
  not NOT_823(g6149,I10810);
  not NOT_824(g3988,g3097);
  not NOT_825(I6686,g2246);
  not NOT_826(g6349,I11374);
  not NOT_827(g5674,g5042);
  not NOT_828(g8177,I14410);
  not NOT_829(g3693,g2424);
  not NOT_830(I11034,g5644);
  not NOT_831(g9223,I15943);
  not NOT_832(I14163,g7533);
  not NOT_833(g2291,I6057);
  not NOT_834(I14012,g7438);
  not NOT_835(I11641,g5918);
  not NOT_836(g6848,I12415);
  not NOT_837(I15580,g8985);
  not NOT_838(I13797,g7502);
  not NOT_839(I12331,g6704);
  not NOT_840(g5541,g4814);
  not NOT_841(g3548,g2185);
  not NOT_842(g1684,g1);
  not NOT_843(g1745,g746);
  not NOT_844(g6198,g5335);
  not NOT_845(g1639,g1207);
  not NOT_846(g2344,I6148);
  not NOT_847(g6855,I12436);
  not NOT_848(g6398,I11515);
  not NOT_849(I10541,g5256);
  not NOT_850(I6121,g321);
  not NOT_851(g7263,I13231);
  not NOT_852(g2207,I5920);
  not NOT_853(g5153,I9585);
  not NOT_854(g5680,g5101);
  not NOT_855(I12897,g6962);
  not NOT_856(I12448,g6569);
  not NOT_857(I12961,g6921);
  not NOT_858(I9515,g4301);
  not NOT_859(I9630,g4867);
  not NOT_860(I14789,g8544);
  not NOT_861(g2259,g1325);
  not NOT_862(g9115,I15735);
  not NOT_863(g4014,I7769);
  not NOT_864(I7079,g2532);
  not NOT_865(I12505,g6612);
  not NOT_866(g9315,I16061);
  not NOT_867(g1808,g629);
  not NOT_868(g4885,g4070);
  not NOT_869(I13635,g7243);
  not NOT_870(g5744,I10289);
  not NOT_871(g8199,I14424);
  not NOT_872(g9047,I15543);
  not NOT_873(g5802,I10445);
  not NOT_874(g4660,I8895);
  not NOT_875(g2923,I6657);
  not NOT_876(I12717,g6543);
  not NOT_877(g1707,g955);
  not NOT_878(I14325,g7713);
  not NOT_879(I10829,g5224);
  not NOT_880(g8781,g8585);
  not NOT_881(I10535,g5254);
  not NOT_882(I5389,g690);
  not NOT_883(I5706,g901);
  not NOT_884(g8898,I15308);
  not NOT_885(g4903,g4084);
  not NOT_886(g7562,I13858);
  not NOT_887(I15178,g8753);
  not NOT_888(I10946,g5563);
  not NOT_889(g8797,I15003);
  not NOT_890(g6524,I11710);
  not NOT_891(I14828,g8639);
  not NOT_892(g6644,g6208);
  not NOT_893(g8510,I14643);
  not NOT_894(I13164,g7086);
  not NOT_895(I5371,g633);
  not NOT_896(g7723,I14042);
  not NOT_897(I14121,g7587);
  not NOT_898(g2215,g1416);
  not NOT_899(I15953,g9215);
  not NOT_900(g6319,I11284);
  not NOT_901(g7101,I12891);
  not NOT_902(g2886,g2240);
  not NOT_903(g3908,I7517);
  not NOT_904(g7301,I13335);
  not NOT_905(I7356,g2843);
  not NOT_906(I13891,g7336);
  not NOT_907(I15654,g9057);
  not NOT_908(g4036,g3192);
  not NOT_909(g6152,I10815);
  not NOT_910(g6258,g5427);
  not NOT_911(g6352,I11383);
  not NOT_912(g6818,I12325);
  not NOT_913(g1575,g685);
  not NOT_914(g1865,g1013);
  not NOT_915(I8483,g3641);
  not NOT_916(g6867,I12472);
  not NOT_917(g3567,g2407);
  not NOT_918(I15417,g8893);
  not NOT_919(g1715,I5559);
  not NOT_920(g2314,I6099);
  not NOT_921(I9440,g4285);
  not NOT_922(I14291,g7680);
  not NOT_923(I12433,g6632);
  not NOT_924(g4335,g3659);
  not NOT_925(I9123,g4455);
  not NOT_926(I15334,g8800);
  not NOT_927(g7751,I14124);
  not NOT_928(g2870,g2225);
  not NOT_929(g5492,g4919);
  not NOT_930(I12148,g5988);
  not NOT_931(I13109,g7059);
  not NOT_932(g4382,I8373);
  not NOT_933(g1833,g770);
  not NOT_934(g5600,g5128);
  not NOT_935(I13537,g7152);
  not NOT_936(g5574,g4969);
  not NOT_937(I8790,g4020);
  not NOT_938(g6211,g5645);
  not NOT_939(g2825,I6553);
  not NOT_940(g2650,I6434);
  not NOT_941(g6186,I10919);
  not NOT_942(g6386,I11485);
  not NOT_943(I12646,g6493);
  not NOT_944(g7585,I13900);
  not NOT_945(g9017,I15475);
  not NOT_946(I9666,g4931);
  not NOT_947(I15762,g9039);
  not NOT_948(I12343,g6731);
  not NOT_949(g4805,I9136);
  not NOT_950(g6975,I12712);
  not NOT_951(g4916,g4202);
  not NOT_952(g4022,I7785);
  not NOT_953(g3965,I7676);
  not NOT_954(I5963,g225);
  not NOT_955(g1584,g738);
  not NOT_956(g6599,I11809);
  not NOT_957(g1896,g86);
  not NOT_958(g7441,I13580);
  not NOT_959(I15423,g8894);
  not NOT_960(g6026,g5384);
  not NOT_961(I9528,g4006);
  not NOT_962(g6426,I11559);
  not NOT_963(I6860,g2185);
  not NOT_964(g3264,I6900);
  not NOT_965(I7053,g2452);
  not NOT_966(I6341,g1351);
  not NOT_967(I10506,g5236);
  not NOT_968(g5580,g4938);
  not NOT_969(I9648,g4795);
  not NOT_970(g9234,I15956);
  not NOT_971(I10028,g4825);
  not NOT_972(g9128,I15762);
  not NOT_973(g6614,I11838);
  not NOT_974(g6370,I11437);
  not NOT_975(I14028,g7501);
  not NOT_976(g3933,g3131);
  not NOT_977(I8904,g4126);
  not NOT_978(g9330,g9319);
  not NOT_979(g6325,I11302);
  not NOT_980(g6821,I12334);
  not NOT_981(g3521,g2185);
  not NOT_982(g4560,g2899);
  not NOT_983(I8446,g3014);
  not NOT_984(g3050,I6788);
  not NOT_985(g3641,I7115);
  not NOT_986(I15909,g9201);
  not NOT_987(I15543,g9006);
  not NOT_988(g5736,I10265);
  not NOT_989(g2943,g2362);
  not NOT_990(g6984,I12725);
  not NOT_991(g7168,I13072);
  not NOT_992(g6939,g6543);
  not NOT_993(g3996,I7731);
  not NOT_994(I11796,g6287);
  not NOT_995(I12412,g6404);
  not NOT_996(I8841,g3979);
  not NOT_997(g5623,g4969);
  not NOT_998(g7772,I14187);
  not NOT_999(g6083,I10702);
  not NOT_1000(g7058,g6649);
  not NOT_1001(I5957,g110);
  not NOT_1002(g2887,g2241);
  not NOT_1003(g4873,I9217);
  not NOT_1004(g4632,I8811);
  not NOT_1005(g7531,I13773);
  not NOT_1006(g4095,I7908);
  not NOT_1007(g5076,I9446);
  not NOT_1008(g8870,I15196);
  not NOT_1009(I8763,g3947);
  not NOT_1010(g4037,g2845);
  not NOT_1011(g6483,I11645);
  not NOT_1012(I12229,g6659);
  not NOT_1013(I9884,g4868);
  not NOT_1014(g2934,I6676);
  not NOT_1015(g5476,g4907);
  not NOT_1016(g7743,I14100);
  not NOT_1017(g4653,I8874);
  not NOT_1018(I6358,g13);
  not NOT_1019(g4102,I7919);
  not NOT_1020(g6636,I11900);
  not NOT_1021(I15568,g8981);
  not NOT_1022(I15747,g9042);
  not NOT_1023(I5865,g1206);
  not NOT_1024(g9213,I15915);
  not NOT_1025(g6106,g5345);
  not NOT_1026(g5175,I9651);
  not NOT_1027(g4579,g2918);
  not NOT_1028(I10649,g5657);
  not NOT_1029(I12011,g5939);
  not NOT_1030(g6306,I11245);
  not NOT_1031(I5715,g896);
  not NOT_1032(g7505,I13695);
  not NOT_1033(g5871,I10558);
  not NOT_1034(g3878,g2962);
  not NOT_1035(g8008,g7559);
  not NOT_1036(g4719,I9021);
  not NOT_1037(g6790,I12241);
  not NOT_1038(g7734,I14073);
  not NOT_1039(I6587,g1708);
  not NOT_1040(g3777,g2170);
  not NOT_1041(g7411,g7202);
  not NOT_1042(I9372,g3902);
  not NOT_1043(I10491,g5231);
  not NOT_1044(I15814,g9154);
  not NOT_1045(g3835,I7308);
  not NOT_1046(I16116,g9350);
  not NOT_1047(g6387,I11488);
  not NOT_1048(I11522,g5847);
  not NOT_1049(g2096,g1226);
  not NOT_1050(I9618,g4742);
  not NOT_1051(I12582,g6745);
  not NOT_1052(g5285,g4841);
  not NOT_1053(g6461,I11607);
  not NOT_1054(g8768,g8585);
  not NOT_1055(I13663,g7235);
  not NOT_1056(g3882,g2970);
  not NOT_1057(g2496,g942);
  not NOT_1058(I7626,g3632);
  not NOT_1059(g4917,g4102);
  not NOT_1060(I15974,g9234);
  not NOT_1061(I6615,g1983);
  not NOT_1062(g6756,I12141);
  not NOT_1063(g8972,I15420);
  not NOT_1064(I10770,g5441);
  not NOT_1065(I12310,g6723);
  not NOT_1066(g1897,g789);
  not NOT_1067(g9090,I15660);
  not NOT_1068(g6622,I11858);
  not NOT_1069(g7474,I13628);
  not NOT_1070(I8757,g3921);
  not NOT_1071(g6027,g5384);
  not NOT_1072(g7992,g7557);
  not NOT_1073(g4265,g3591);
  not NOT_1074(g3611,I7079);
  not NOT_1075(g6427,I11562);
  not NOT_1076(g2137,I5889);
  not NOT_1077(g2891,g2265);
  not NOT_1078(g5184,I9678);
  not NOT_1079(I15638,g8978);
  not NOT_1080(g9366,I16126);
  not NOT_1081(g2913,g2307);
  not NOT_1082(I12379,g6768);
  not NOT_1083(g5139,I9543);
  not NOT_1084(g5384,I9837);
  not NOT_1085(g6904,g6426);
  not NOT_1086(I12958,g6920);
  not NOT_1087(g9056,I15562);
  not NOT_1088(g8065,I14338);
  not NOT_1089(I8315,g3691);
  not NOT_1090(I8811,g4022);
  not NOT_1091(g6446,I11591);
  not NOT_1092(g8228,I14463);
  not NOT_1093(g3981,I7706);
  not NOT_1094(g5024,I9360);
  not NOT_1095(g6514,I11696);
  not NOT_1096(I6239,g8);
  not NOT_1097(g3674,I7164);
  not NOT_1098(g2807,g1782);
  not NOT_1099(I5362,g3841);
  not NOT_1100(I11326,g5819);
  not NOT_1101(I9555,g4892);
  not NOT_1102(g5795,I10424);
  not NOT_1103(g5737,I10268);
  not NOT_1104(I15391,g8917);
  not NOT_1105(g6403,I11522);
  not NOT_1106(I13326,g7176);
  not NOT_1107(g5809,I10460);
  not NOT_1108(I5419,g1603);
  not NOT_1109(I9804,g5113);
  not NOT_1110(I10262,g5551);
  not NOT_1111(I7683,g2573);
  not NOT_1112(g3997,I7734);
  not NOT_1113(I12742,g6590);
  not NOT_1114(g6345,I11362);
  not NOT_1115(g6841,I12394);
  not NOT_1116(I15510,g8969);
  not NOT_1117(I11040,g5299);
  not NOT_1118(I11948,g5897);
  not NOT_1119(I8874,g3884);
  not NOT_1120(g2266,I6003);
  not NOT_1121(g6763,I12158);
  not NOT_1122(I7778,g3019);
  not NOT_1123(I16142,g9366);
  not NOT_1124(g6391,I11500);
  not NOT_1125(g1006,I5410);
  not NOT_1126(g4296,g3790);
  not NOT_1127(I6853,g2185);
  not NOT_1128(g3238,I6894);
  not NOT_1129(I9621,g4732);
  not NOT_1130(g5477,g4908);
  not NOT_1131(g9260,I15990);
  not NOT_1132(g5523,I9935);
  not NOT_1133(I12681,g6469);
  not NOT_1134(I10719,g5559);
  not NOT_1135(g6637,I11903);
  not NOT_1136(g5643,I10128);
  not NOT_1137(I15014,g8607);
  not NOT_1138(g1801,g618);
  not NOT_1139(g4553,g2891);
  not NOT_1140(g9063,I15583);
  not NOT_1141(g6307,I11248);
  not NOT_1142(I15586,g8987);
  not NOT_1143(I15007,g8627);
  not NOT_1144(I8880,g4303);
  not NOT_1145(I14718,g8068);
  not NOT_1146(g3802,g1832);
  not NOT_1147(g7688,g7406);
  not NOT_1148(g6359,I11404);
  not NOT_1149(g6223,I11008);
  not NOT_1150(g2481,I6317);
  not NOT_1151(g8913,I15329);
  not NOT_1152(g1748,g601);
  not NOT_1153(g2692,g1671);
  not NOT_1154(g4012,I7765);
  not NOT_1155(g6858,I12445);
  not NOT_1156(g5742,I10283);
  not NOT_1157(g5551,I9974);
  not NOT_1158(g5099,g4477);
  not NOT_1159(g2497,g945);
  not NOT_1160(I12690,g6467);
  not NOT_1161(g2354,I6178);
  not NOT_1162(I16165,g9377);
  not NOT_1163(g2960,g2381);
  not NOT_1164(g4706,I9005);
  not NOT_1165(I9567,g4693);
  not NOT_1166(I7526,g2752);
  not NOT_1167(I5897,g173);
  not NOT_1168(I14573,g8179);
  not NOT_1169(I10247,g5266);
  not NOT_1170(g3901,I7492);
  not NOT_1171(g7000,I12742);
  not NOT_1172(I13509,g7137);
  not NOT_1173(I15720,g9053);
  not NOT_1174(g9318,g9304);
  not NOT_1175(g9367,I16129);
  not NOT_1176(I11933,g5847);
  not NOT_1177(g7126,I12968);
  not NOT_1178(I8935,g4005);
  not NOT_1179(I5425,g1245);
  not NOT_1180(g4029,I7800);
  not NOT_1181(g6251,I11060);
  not NOT_1182(g6315,I11272);
  not NOT_1183(g6811,I12304);
  not NOT_1184(g6642,I11912);
  not NOT_1185(g4371,I8354);
  not NOT_1186(I11851,g6277);
  not NOT_1187(g3511,g1616);
  not NOT_1188(g5754,g5403);
  not NOT_1189(g9057,I15565);
  not NOT_1190(I16006,g9261);
  not NOT_1191(g7760,I14151);
  not NOT_1192(I14388,g7605);
  not NOT_1193(I7850,g2795);
  not NOT_1194(g9193,g9181);
  not NOT_1195(g3092,I6826);
  not NOT_1196(I14777,g8511);
  not NOT_1197(g3492,I6970);
  not NOT_1198(g4281,g2562);
  not NOT_1199(g6874,I12493);
  not NOT_1200(g5613,g4748);
  not NOT_1201(I14251,g7541);
  not NOT_1202(g3574,g1771);
  not NOT_1203(g3864,g2943);
  not NOT_1204(g8342,g8008);
  not NOT_1205(I15340,g8856);
  not NOT_1206(g2267,I6006);
  not NOT_1207(g2312,I6093);
  not NOT_1208(g6654,I11942);
  not NOT_1209(g5444,g5074);
  not NOT_1210(g5269,I9791);
  not NOT_1211(I7702,g3062);
  not NOT_1212(I15684,g9067);
  not NOT_1213(g8481,I14637);
  not NOT_1214(I12128,g5897);
  not NOT_1215(g1578,g699);
  not NOT_1216(g1868,I5747);
  not NOT_1217(I9360,g4257);
  not NOT_1218(g2401,g22);
  not NOT_1219(I7919,g3761);
  not NOT_1220(I10032,g1236);
  not NOT_1221(g1718,I5562);
  not NOT_1222(g7779,I14208);
  not NOT_1223(g2293,g888);
  not NOT_1224(g6880,I12511);
  not NOT_1225(g4684,I8949);
  not NOT_1226(I9050,g3881);
  not NOT_1227(I11452,g6071);
  not NOT_1228(g6595,g6083);
  not NOT_1229(g4639,I8832);
  not NOT_1230(I5682,g168);
  not NOT_1231(I5766,g1254);
  not NOT_1232(I11047,g5653);
  not NOT_1233(I13574,g7205);
  not NOT_1234(g2329,I6130);
  not NOT_1235(I6440,g1806);
  not NOT_1236(g7023,I12779);
  not NOT_1237(g9121,I15747);
  not NOT_1238(g4963,g4328);
  not NOT_1239(g2761,g1820);
  not NOT_1240(I5801,g1424);
  not NOT_1241(g9321,g9311);
  not NOT_1242(g8960,I15394);
  not NOT_1243(g7423,I13544);
  not NOT_1244(g1582,g714);
  not NOT_1245(I11912,g5897);
  not NOT_1246(I11311,g5760);
  not NOT_1247(I13912,g7359);
  not NOT_1248(I13311,g7162);
  not NOT_1249(g2828,g1980);
  not NOT_1250(I12298,g6697);
  not NOT_1251(I6323,g1342);
  not NOT_1252(I14061,g7546);
  not NOT_1253(g1793,g626);
  not NOT_1254(I7561,g2562);
  not NOT_1255(g7588,I13909);
  not NOT_1256(I10766,g5674);
  not NOT_1257(g2727,g2424);
  not NOT_1258(g4808,I9145);
  not NOT_1259(g6978,I12717);
  not NOT_1260(g6612,I11832);
  not NOT_1261(g7161,I13057);
  not NOT_1262(g1015,I5416);
  not NOT_1263(g5729,g5144);
  not NOT_1264(g3968,I7683);
  not NOT_1265(g6243,I11050);
  not NOT_1266(g7361,I13499);
  not NOT_1267(I15193,g8774);
  not NOT_1268(I13051,g6967);
  not NOT_1269(I13072,g6969);
  not NOT_1270(g2746,g2259);
  not NOT_1271(I12737,g6460);
  not NOT_1272(g2221,I5936);
  not NOT_1273(g3076,g1831);
  not NOT_1274(g7127,g6974);
  not NOT_1275(g8783,g8524);
  not NOT_1276(g7327,I13403);
  not NOT_1277(I12232,g6662);
  not NOT_1278(g1664,g1462);
  not NOT_1279(I6151,g12);
  not NOT_1280(g1246,I5425);
  not NOT_1281(g2703,g1809);
  not NOT_1282(g8218,I14433);
  not NOT_1283(I8823,g3965);
  not NOT_1284(g5014,I9344);
  not NOT_1285(g206,I5353);
  not NOT_1286(g6328,I11311);
  not NOT_1287(g6130,I10761);
  not NOT_1288(g7146,g6998);
  not NOT_1289(g6542,I11718);
  not NOT_1290(g6330,I11317);
  not NOT_1291(g7346,I13454);
  not NOT_1292(g7633,I13962);
  not NOT_1293(g1721,I5565);
  not NOT_1294(I11350,g5763);
  not NOT_1295(g3871,g2953);
  not NOT_1296(I7970,g3557);
  not NOT_1297(I13350,g7223);
  not NOT_1298(I15475,g8901);
  not NOT_1299(g2932,g2329);
  not NOT_1300(g7103,I12897);
  not NOT_1301(I9271,g4263);
  not NOT_1302(g3651,I7129);
  not NOT_1303(g7303,I13341);
  not NOT_1304(I7925,g2761);
  not NOT_1305(g8676,I14822);
  not NOT_1306(g2624,g1569);
  not NOT_1307(g2953,g2373);
  not NOT_1308(I15222,g8834);
  not NOT_1309(g6800,I12271);
  not NOT_1310(g3285,g1689);
  not NOT_1311(I13152,g6966);
  not NOT_1312(g8761,g8564);
  not NOT_1313(g4604,I8727);
  not NOT_1314(I10451,g5216);
  not NOT_1315(I10472,g5223);
  not NOT_1316(I13846,g7487);
  not NOT_1317(g3500,g1616);
  not NOT_1318(I14451,g8172);
  not NOT_1319(g7732,I14067);
  not NOT_1320(I5407,g4653);
  not NOT_1321(I13731,g7441);
  not NOT_1322(I5920,g219);
  not NOT_1323(I6839,g2185);
  not NOT_1324(I5868,g74);
  not NOT_1325(I7320,g2927);
  not NOT_1326(g2677,g1664);
  not NOT_1327(g7753,I14130);
  not NOT_1328(g5178,I9660);
  not NOT_1329(g5679,I10172);
  not NOT_1330(I11413,g5871);
  not NOT_1331(I5718,g896);
  not NOT_1332(g7508,I13704);
  not NOT_1333(I13413,g7127);
  not NOT_1334(g6213,I10976);
  not NOT_1335(I5535,g48);
  not NOT_1336(g2866,g2221);
  not NOT_1337(g4584,g3466);
  not NOT_1338(I12445,g6568);
  not NOT_1339(g4539,g2881);
  not NOT_1340(g8746,g8524);
  not NOT_1341(g8221,I14442);
  not NOT_1342(g5335,g4677);
  not NOT_1343(g5831,I10516);
  not NOT_1344(g3838,I7317);
  not NOT_1345(g1689,g855);
  not NOT_1346(g2149,I5894);
  not NOT_1347(g2349,I6163);
  not NOT_1348(I12499,g6597);
  not NOT_1349(g7043,g6543);
  not NOT_1350(g9141,g9129);
  not NOT_1351(g5182,I9672);
  not NOT_1352(I10776,g5576);
  not NOT_1353(I12316,g6736);
  not NOT_1354(I9132,g4284);
  not NOT_1355(I6143,g1217);
  not NOT_1356(I9209,g4349);
  not NOT_1357(g7116,I12936);
  not NOT_1358(g1671,g1494);
  not NOT_1359(I7987,g3528);
  not NOT_1360(g5805,I10448);
  not NOT_1361(g5916,g5384);
  not NOT_1362(g5022,g4438);
  not NOT_1363(g2699,g1674);
  not NOT_1364(g4019,I7778);
  not NOT_1365(g6090,g5529);
  not NOT_1366(g4362,g2810);
  not NOT_1367(I11929,g6190);
  not NOT_1368(I12989,g6932);
  not NOT_1369(g3077,I6805);
  not NOT_1370(g7034,g6525);
  not NOT_1371(g5749,g5207);
  not NOT_1372(g6490,I11656);
  not NOT_1373(g6823,I12340);
  not NOT_1374(g7434,I13565);
  not NOT_1375(I14825,g8651);
  not NOT_1376(g3523,g2407);
  not NOT_1377(I14370,g7603);
  not NOT_1378(g6366,I11425);
  not NOT_1379(I12722,g6611);
  not NOT_1380(g7565,I13865);
  not NOT_1381(I7299,g2961);
  not NOT_1382(I5664,g916);
  not NOT_1383(g3643,g2453);
  not NOT_1384(I12924,g6983);
  not NOT_1385(I13583,g7252);
  not NOT_1386(g2241,I5984);
  not NOT_1387(g1564,g642);
  not NOT_1388(g7147,g6904);
  not NOT_1389(I16122,g9353);
  not NOT_1390(I10151,g5007);
  not NOT_1391(I10172,g4873);
  not NOT_1392(g7347,I13457);
  not NOT_1393(I15516,g8977);
  not NOT_1394(I9558,g4597);
  not NOT_1395(g5798,I10433);
  not NOT_1396(I14151,g7555);
  not NOT_1397(g1826,g632);
  not NOT_1398(I12271,g6663);
  not NOT_1399(I14172,g7545);
  not NOT_1400(g6148,I10807);
  not NOT_1401(g6649,I11929);
  not NOT_1402(I14996,g8510);
  not NOT_1403(g6348,I11371);
  not NOT_1404(I8989,g4537);
  not NOT_1405(g8677,I14825);
  not NOT_1406(g7533,I13779);
  not NOT_1407(g3634,I7107);
  not NOT_1408(I8193,g3547);
  not NOT_1409(g6155,I10826);
  not NOT_1410(I14844,g8641);
  not NOT_1411(g6851,I12424);
  not NOT_1412(g6355,I11392);
  not NOT_1413(I11787,g6273);
  not NOT_1414(I14394,g7536);
  not NOT_1415(I12753,g6445);
  not NOT_1416(g8866,I15184);
  not NOT_1417(g7210,I13144);
  not NOT_1418(g2644,I6416);
  not NOT_1419(g3499,g2185);
  not NOT_1420(I8971,g4464);
  not NOT_1421(I12145,g5971);
  not NOT_1422(g1638,g1092);
  not NOT_1423(I11302,g5796);
  not NOT_1424(I7738,g3038);
  not NOT_1425(g5873,g5367);
  not NOT_1426(I13302,g7164);
  not NOT_1427(g5037,g4438);
  not NOT_1428(g9111,I15723);
  not NOT_1429(I12199,g6475);
  not NOT_1430(g7013,I12757);
  not NOT_1431(g9311,I16049);
  not NOT_1432(g5437,g5041);
  not NOT_1433(I11827,g6231);
  not NOT_1434(g5653,g4748);
  not NOT_1435(g7413,I13524);
  not NOT_1436(I13743,g7454);
  not NOT_1437(g3926,I7581);
  not NOT_1438(g5302,g5028);
  not NOT_1439(I14420,g7554);
  not NOT_1440(I15208,g8810);
  not NOT_1441(g2818,g1792);
  not NOT_1442(g6063,I10678);
  not NOT_1443(g4070,I7847);
  not NOT_1444(I12529,g6628);
  not NOT_1445(g2867,g2222);
  not NOT_1446(g3754,g2543);
  not NOT_1447(I9600,g4698);
  not NOT_1448(g8198,g7721);
  not NOT_1449(g8747,g8545);
  not NOT_1450(g4025,I7792);
  not NOT_1451(I14318,g7657);
  not NOT_1452(g5719,I10236);
  not NOT_1453(I12696,g6503);
  not NOT_1454(g9374,I16148);
  not NOT_1455(I14227,g7552);
  not NOT_1456(I5689,g906);
  not NOT_1457(I7959,g2793);
  not NOT_1458(g1758,g1084);
  not NOT_1459(g1589,g746);
  not NOT_1460(I14025,g7500);
  not NOT_1461(I7517,g3578);
  not NOT_1462(I11803,g6280);
  not NOT_1463(I7082,g2470);
  not NOT_1464(g2893,I6615);
  not NOT_1465(I15726,g9069);
  not NOT_1466(g7117,I12939);
  not NOT_1467(g6279,I11132);
  not NOT_1468(g5917,g5412);
  not NOT_1469(g7317,I13383);
  not NOT_1470(I14058,g7544);
  not NOT_1471(g6720,g6254);
  not NOT_1472(I5428,g49);
  not NOT_1473(g6118,g5549);
  not NOT_1474(g6167,I10862);
  not NOT_1475(g6318,I11281);
  not NOT_1476(g1571,g669);
  not NOT_1477(g3983,g2845);
  not NOT_1478(g6367,I11428);
  not NOT_1479(g9180,I15824);
  not NOT_1480(g6872,I12487);
  not NOT_1481(g7601,g7450);
  not NOT_1482(I15607,g8994);
  not NOT_1483(g9380,g9379);
  not NOT_1484(g3862,I7389);
  not NOT_1485(g5042,I9396);
  not NOT_1486(g1711,I5555);
  not NOT_1487(g2274,g782);
  not NOT_1488(g6652,I11936);
  not NOT_1489(I12161,g5971);
  not NOT_1490(g4678,I8935);
  not NOT_1491(g3712,g1952);
  not NOT_1492(g8524,g7855);
  not NOT_1493(g6843,I12400);
  not NOT_1494(I15530,g8972);
  not NOT_1495(g5786,I10403);
  not NOT_1496(g4006,I7749);
  not NOT_1497(g2170,g1229);
  not NOT_1498(g1827,g762);
  not NOT_1499(g2614,g1562);
  not NOT_1500(g9020,I15484);
  not NOT_1501(g7775,I14196);
  not NOT_1502(g5164,I9618);
  not NOT_1503(g6393,I11506);
  not NOT_1504(g4635,I8820);
  not NOT_1505(g5364,g5124);
  not NOT_1506(I15565,g8980);
  not NOT_1507(g2325,I6118);
  not NOT_1508(g2821,g1786);
  not NOT_1509(I12259,g6652);
  not NOT_1510(I10377,g5188);
  not NOT_1511(g1774,I5616);
  not NOT_1512(I12708,g6482);
  not NOT_1513(g7581,I13888);
  not NOT_1514(I11662,g5956);
  not NOT_1515(I10739,g5572);
  not NOT_1516(g4087,I7882);
  not NOT_1517(g4105,I7928);
  not NOT_1518(g8152,I14388);
  not NOT_1519(I9076,g4353);
  not NOT_1520(g5054,g4457);
  not NOT_1521(g6834,I12373);
  not NOT_1522(g4801,I9126);
  not NOT_1523(g8867,I15187);
  not NOT_1524(I9889,g4819);
  not NOT_1525(I14739,g8173);
  not NOT_1526(g2939,g2348);
  not NOT_1527(g3961,g3131);
  not NOT_1528(g7060,g6654);
  not NOT_1529(I11890,g6135);
  not NOT_1530(g1803,g758);
  not NOT_1531(g7460,g7172);
  not NOT_1532(I15641,g9017);
  not NOT_1533(I6160,g324);
  not NOT_1534(g5725,g4841);
  not NOT_1535(g4748,g4465);
  not NOT_1536(I11482,g6117);
  not NOT_1537(g6598,I11806);
  not NOT_1538(g3927,I7584);
  not NOT_1539(I5609,g16);
  not NOT_1540(I11248,g6149);
  not NOT_1541(g1780,g614);
  not NOT_1542(I12244,g6642);
  not NOT_1543(I11710,g6098);
  not NOT_1544(I13710,g7340);
  not NOT_1545(g2636,g1580);
  not NOT_1546(g7739,I14088);
  not NOT_1547(g3014,I6767);
  not NOT_1548(I9651,g4805);
  not NOT_1549(g6321,I11290);
  not NOT_1550(g4226,g3591);
  not NOT_1551(g8386,g8014);
  not NOT_1552(I5883,g80);
  not NOT_1553(g2106,I5883);
  not NOT_1554(g8975,I15429);
  not NOT_1555(g3946,g3097);
  not NOT_1556(g2306,I6075);
  not NOT_1557(I13779,g7406);
  not NOT_1558(g9204,I15894);
  not NOT_1559(I15408,g8896);
  not NOT_1560(I15635,g8976);
  not NOT_1561(g6625,I11867);
  not NOT_1562(g1662,g1412);
  not NOT_1563(g2790,g1793);
  not NOT_1564(g7937,I14285);
  not NOT_1565(I7762,g3029);
  not NOT_1566(I12810,g6607);
  not NOT_1567(g6232,I11031);
  not NOT_1568(I11778,g6180);
  not NOT_1569(g3903,I7498);
  not NOT_1570(g9100,I15690);
  not NOT_1571(I12068,g5847);
  not NOT_1572(I10427,g5210);
  not NOT_1573(g7479,I13635);
  not NOT_1574(g9300,I16026);
  not NOT_1575(g5412,I9850);
  not NOT_1576(I10366,g5715);
  not NOT_1577(g6253,g5403);
  not NOT_1578(g6938,I12635);
  not NOT_1579(I14427,g7835);
  not NOT_1580(I5466,g926);
  not NOT_1581(g6813,I12310);
  not NOT_1582(g7294,I13314);
  not NOT_1583(g4373,I8360);
  not NOT_1584(g3513,g2407);
  not NOT_1585(I9139,g4364);
  not NOT_1586(g6909,I12592);
  not NOT_1587(g7190,I13112);
  not NOT_1588(g2622,g1568);
  not NOT_1589(I11945,g5874);
  not NOT_1590(I12337,g6724);
  not NOT_1591(I5365,g3843);
  not NOT_1592(I5861,g1313);
  not NOT_1593(I11356,g5799);
  not NOT_1594(I13356,g7221);
  not NOT_1595(g1816,g767);
  not NOT_1596(g5171,I9639);
  not NOT_1597(g4602,I8721);
  not NOT_1598(g7501,I13679);
  not NOT_1599(I11380,g5822);
  not NOT_1600(I10403,g5202);
  not NOT_1601(g5787,I10406);
  not NOT_1602(g4007,I7752);
  not NOT_1603(g2904,g2287);
  not NOT_1604(I14403,g7679);
  not NOT_1605(g7156,I13042);
  not NOT_1606(g5956,I10582);
  not NOT_1607(g6552,I11722);
  not NOT_1608(g7356,I13484);
  not NOT_1609(g4920,g4105);
  not NOT_1610(g6606,I11824);
  not NOT_1611(g4578,g2917);
  not NOT_1612(I11090,g1000);
  not NOT_1613(I7928,g2873);
  not NOT_1614(I11998,g5918);
  not NOT_1615(g8544,I14657);
  not NOT_1616(g3831,I7296);
  not NOT_1617(I11233,g6147);
  not NOT_1618(g2514,g1330);
  not NOT_1619(g4718,I9018);
  not NOT_1620(g8483,g8038);
  not NOT_1621(I8962,g4553);
  not NOT_1622(I7064,g2458);
  not NOT_1623(I11672,g5971);
  not NOT_1624(g1847,g765);
  not NOT_1625(I9672,g4803);
  not NOT_1626(I15711,g9075);
  not NOT_1627(I13672,g7242);
  not NOT_1628(I7899,g3743);
  not NOT_1629(g4535,g2876);
  not NOT_1630(g2403,g1176);
  not NOT_1631(g8636,I14718);
  not NOT_1632(g1685,I5528);
  not NOT_1633(g2145,g1296);
  not NOT_1634(g6687,I12003);
  not NOT_1635(g2345,I6151);
  not NOT_1636(g2841,g2208);
  not NOT_1637(I7785,g3029);
  not NOT_1638(g7704,I14001);
  not NOT_1639(g4582,g2922);
  not NOT_1640(g3805,g1752);
  not NOT_1641(g3916,I7545);
  not NOT_1642(g9323,g9315);
  not NOT_1643(g6586,I11778);
  not NOT_1644(g8790,g8585);
  not NOT_1645(g2695,g1672);
  not NOT_1646(g4015,g3160);
  not NOT_1647(g2637,g1581);
  not NOT_1648(I11449,g6068);
  not NOT_1649(I12918,g7013);
  not NOT_1650(g5684,I10183);
  not NOT_1651(g8061,I14330);
  not NOT_1652(g5745,I10292);
  not NOT_1653(I15492,g8971);
  not NOT_1654(g5639,g4748);
  not NOT_1655(I14127,g7594);
  not NOT_1656(g7163,I13063);
  not NOT_1657(g3947,I7640);
  not NOT_1658(I11897,g6141);
  not NOT_1659(g2307,I6078);
  not NOT_1660(I11961,g5988);
  not NOT_1661(g7032,g6525);
  not NOT_1662(g2536,g1354);
  not NOT_1663(g5109,I9493);
  not NOT_1664(I13897,g7354);
  not NOT_1665(g8756,g8564);
  not NOT_1666(g3798,g1757);
  not NOT_1667(g5309,g4969);
  not NOT_1668(g7432,I13559);
  not NOT_1669(g6141,I10786);
  not NOT_1670(g6860,I12451);
  not NOT_1671(g2359,g1397);
  not NOT_1672(g4664,I8907);
  not NOT_1673(I9499,g4382);
  not NOT_1674(g6341,I11350);
  not NOT_1675(I11404,g5834);
  not NOT_1676(g3560,g2361);
  not NOT_1677(g9351,I16103);
  not NOT_1678(g2223,I5942);
  not NOT_1679(I7844,g3784);
  not NOT_1680(I15982,g9236);
  not NOT_1681(g5808,I10457);
  not NOT_1682(g1562,g636);
  not NOT_1683(I6680,g1558);
  not NOT_1684(g6645,I11917);
  not NOT_1685(I16040,g9285);
  not NOT_1686(g4721,I9025);
  not NOT_1687(I14103,g7584);
  not NOT_1688(I11212,g6146);
  not NOT_1689(g2016,I5852);
  not NOT_1690(I7731,g3029);
  not NOT_1691(g5759,I10350);
  not NOT_1692(g8514,g8040);
  not NOT_1693(g3873,g2956);
  not NOT_1694(g3632,I7101);
  not NOT_1695(g3095,I6831);
  not NOT_1696(g1817,I5689);
  not NOT_1697(g3495,g1616);
  not NOT_1698(g3653,g2459);
  not NOT_1699(I8180,g3529);
  not NOT_1700(I12322,g6751);
  not NOT_1701(g8145,I14381);
  not NOT_1702(g2522,g1342);
  not NOT_1703(I14181,g7725);
  not NOT_1704(g7157,I13045);
  not NOT_1705(g2642,g1588);
  not NOT_1706(I8832,g3936);
  not NOT_1707(g6879,I12508);
  not NOT_1708(g7357,I13487);
  not NOT_1709(g6607,I11827);
  not NOT_1710(I12532,g6594);
  not NOT_1711(g3579,g1929);
  not NOT_1712(g3869,I7400);
  not NOT_1713(g6962,I12687);
  not NOT_1714(I8853,g4034);
  not NOT_1715(g6659,I11955);
  not NOT_1716(I12158,g5956);
  not NOT_1717(g6358,I11401);
  not NOT_1718(g6506,I11680);
  not NOT_1719(g1751,g452);
  not NOT_1720(I5847,g1360);
  not NOT_1721(I12561,g6449);
  not NOT_1722(I16183,g9388);
  not NOT_1723(g5604,g4969);
  not NOT_1724(I12295,g6693);
  not NOT_1725(g3917,I7548);
  not NOT_1726(g2654,I6446);
  not NOT_1727(I10190,g4670);
  not NOT_1728(g1585,g724);
  not NOT_1729(g4689,I8966);
  not NOT_1730(g6587,I11781);
  not NOT_1731(g9372,I16142);
  not NOT_1732(I15522,g9018);
  not NOT_1733(I15663,g9066);
  not NOT_1734(I14190,g7531);
  not NOT_1735(I9543,g4279);
  not NOT_1736(g6111,g5453);
  not NOT_1737(g8223,I14448);
  not NOT_1738(g6311,I11260);
  not NOT_1739(g5833,I10522);
  not NOT_1740(I7814,g2605);
  not NOT_1741(I13646,g7245);
  not NOT_1742(g9235,I15959);
  not NOT_1743(g4028,I7797);
  not NOT_1744(g2880,g2234);
  not NOT_1745(I7350,g2971);
  not NOT_1746(I6574,g576);
  not NOT_1747(g2595,g1643);
  not NOT_1748(I6864,g2528);
  not NOT_1749(I11971,g6179);
  not NOT_1750(g4030,g3160);
  not NOT_1751(g8016,I14311);
  not NOT_1752(g8757,g8585);
  not NOT_1753(g5584,g4841);
  not NOT_1754(g1673,g1504);
  not NOT_1755(g6374,I11449);
  not NOT_1756(I14211,g7712);
  not NOT_1757(g9134,I15776);
  not NOT_1758(I15553,g9009);
  not NOT_1759(I13369,g7268);
  not NOT_1760(g2272,I6021);
  not NOT_1761(I14088,g7585);
  not NOT_1762(g4564,I8665);
  not NOT_1763(I11368,g5833);
  not NOT_1764(g8642,I14732);
  not NOT_1765(I5562,g1300);
  not NOT_1766(I12364,g6714);
  not NOT_1767(I7769,g3038);
  not NOT_1768(g5162,I9612);
  not NOT_1769(g3770,g2551);
  not NOT_1770(g5268,I9788);
  not NOT_1771(I9014,g3864);
  not NOT_1772(g5362,I9823);
  not NOT_1773(I10497,g5233);
  not NOT_1774(I15536,g9004);
  not NOT_1775(g1772,g607);
  not NOT_1776(g6380,I11467);
  not NOT_1777(I9660,g4806);
  not NOT_1778(g6591,I11787);
  not NOT_1779(I15702,g9064);
  not NOT_1780(I13850,g7328);
  not NOT_1781(g6832,I12367);
  not NOT_1782(I5817,g1081);
  not NOT_1783(g2982,g1848);
  not NOT_1784(g8874,I15208);
  not NOT_1785(g3532,g2407);
  not NOT_1786(I7967,g2787);
  not NOT_1787(g7778,I14205);
  not NOT_1788(g1743,g598);
  not NOT_1789(g2234,I5963);
  not NOT_1790(g6853,I12430);
  not NOT_1791(g2128,g1284);
  not NOT_1792(g4638,I8829);
  not NOT_1793(g2629,g1574);
  not NOT_1794(g6020,g5367);
  not NOT_1795(g2328,I6127);
  not NOT_1796(I10987,g5609);
  not NOT_1797(I12289,g6702);
  not NOT_1798(I5605,g58);
  not NOT_1799(I10250,g5268);
  not NOT_1800(g7735,I14076);
  not NOT_1801(g4609,I8742);
  not NOT_1802(g6507,I11683);
  not NOT_1803(g4308,I8277);
  not NOT_1804(g1011,I5413);
  not NOT_1805(I13228,g6892);
  not NOT_1806(g9113,I15729);
  not NOT_1807(g6794,I12253);
  not NOT_1808(g1856,g774);
  not NOT_1809(I12571,g6729);
  not NOT_1810(g9313,I16055);
  not NOT_1811(I11011,g5693);
  not NOT_1812(I5751,g963);
  not NOT_1813(g5086,I9460);
  not NOT_1814(g8880,I15218);
  not NOT_1815(g3189,I6864);
  not NOT_1816(I13716,g7331);
  not NOT_1817(g5730,I10247);
  not NOT_1818(g7475,I13631);
  not NOT_1819(I16072,g9303);
  not NOT_1820(g3990,g3160);
  not NOT_1821(g2554,I6376);
  not NOT_1822(I14338,g7581);
  not NOT_1823(g5185,I9681);
  not NOT_1824(g4589,g2930);
  not NOT_1825(I10969,g5606);
  not NOT_1826(g9094,I15672);
  not NOT_1827(g7627,I13956);
  not NOT_1828(g3888,g3097);
  not NOT_1829(I15062,g8632);
  not NOT_1830(g6905,I12586);
  not NOT_1831(g3029,g1929);
  not NOT_1832(g7292,I13308);
  not NOT_1833(g3787,g1842);
  not NOT_1834(g8017,g7692);
  not NOT_1835(g6628,I11880);
  not NOT_1836(I15933,g9210);
  not NOT_1837(g7526,I13758);
  not NOT_1838(g5470,g4899);
  not NOT_1839(g5897,I10569);
  not NOT_1840(g3956,g2845);
  not NOT_1841(g5025,I9363);
  not NOT_1842(g6515,g6125);
  not NOT_1843(I11627,g5874);
  not NOT_1844(g6630,I11884);
  not NOT_1845(g4571,g2908);
  not NOT_1846(I12687,g6745);
  not NOT_1847(g3675,I7167);
  not NOT_1848(I12976,g6928);
  not NOT_1849(g1573,g677);
  not NOT_1850(g1863,g68);
  not NOT_1851(g6300,I11227);
  not NOT_1852(I13112,g7021);
  not NOT_1853(g7603,I13940);
  not NOT_1854(I11050,g5335);
  not NOT_1855(I11958,g5874);
  not NOT_1856(g7039,g6543);
  not NOT_1857(I9422,g4360);
  not NOT_1858(I8351,g1160);
  not NOT_1859(g8234,I14489);
  not NOT_1860(g4455,g3811);
  not NOT_1861(g2902,g2285);
  not NOT_1862(g7439,I13574);
  not NOT_1863(I12643,g6501);
  not NOT_1864(I5368,g3853);
  not NOT_1865(I11386,g5764);
  not NOT_1866(g1569,g661);
  not NOT_1867(g453,I5362);
  not NOT_1868(I5772,g1240);
  not NOT_1869(g2490,I6326);
  not NOT_1870(I6024,g544);
  not NOT_1871(I5531,g866);
  not NOT_1872(g2366,I6198);
  not NOT_1873(I12669,g6477);
  not NOT_1874(g7583,I13894);
  not NOT_1875(g7702,I13997);
  not NOT_1876(g4196,I8097);
  not NOT_1877(g5678,I10169);
  not NOT_1878(I6795,g1683);
  not NOT_1879(I10503,g5235);
  not NOT_1880(g3684,g2180);
  not NOT_1881(g3639,g2424);
  not NOT_1882(g4803,I9132);
  not NOT_1883(g6973,I12708);
  not NOT_1884(g5006,I9333);
  not NOT_1885(g3338,g1901);
  not NOT_1886(g8800,I15010);
  not NOT_1887(g3963,I7672);
  not NOT_1888(g9360,I16116);
  not NOT_1889(I15574,g8983);
  not NOT_1890(g4538,g2880);
  not NOT_1891(g1688,I5535);
  not NOT_1892(g2148,g1304);
  not NOT_1893(I15205,g8809);
  not NOT_1894(g2649,I6431);
  not NOT_1895(g4780,I9089);
  not NOT_1896(g1857,g889);
  not NOT_1897(g2348,I6160);
  not NOT_1898(I7788,g2595);
  not NOT_1899(g9050,I15550);
  not NOT_1900(g5682,I10177);
  not NOT_1901(g5766,I10373);
  not NOT_1902(g5087,I9463);
  not NOT_1903(g1976,g1269);
  not NOT_1904(g6969,I12702);
  not NOT_1905(I15912,g9193);
  not NOT_1906(I9095,g4283);
  not NOT_1907(g5801,I10442);
  not NOT_1908(g3808,g1827);
  not NOT_1909(g7276,I13264);
  not NOT_1910(g5487,I9907);
  not NOT_1911(I14315,g7676);
  not NOT_1912(I6643,g1970);
  not NOT_1913(I11793,g6188);
  not NOT_1914(I11428,g5813);
  not NOT_1915(I12424,g6446);
  not NOT_1916(I13428,g7167);
  not NOT_1917(g3707,g2226);
  not NOT_1918(g6323,I11296);
  not NOT_1919(I14819,g8647);
  not NOT_1920(g4662,I8901);
  not NOT_1921(g2698,g1673);
  not NOT_1922(g4018,I7775);
  not NOT_1923(I12558,g6449);
  not NOT_1924(I14202,g7708);
  not NOT_1925(I8172,g3524);
  not NOT_1926(I14257,g7716);
  not NOT_1927(I9579,g4713);
  not NOT_1928(g2964,I6716);
  not NOT_1929(I14055,g7495);
  not NOT_1930(I16020,g9264);
  not NOT_1931(g9379,I16161);
  not NOT_1932(I7392,g3230);
  not NOT_1933(g5755,g5494);
  not NOT_1934(I15592,g8989);
  not NOT_1935(I15756,g9081);
  not NOT_1936(g7527,I13761);
  not NOT_1937(I14070,g7714);
  not NOT_1938(g3957,I7662);
  not NOT_1939(I12544,g6617);
  not NOT_1940(I6099,g584);
  not NOT_1941(I9752,g4705);
  not NOT_1942(g4093,I7902);
  not NOT_1943(g8512,g8094);
  not NOT_1944(I8282,g3515);
  not NOT_1945(I16046,g9288);
  not NOT_1946(g1760,I5605);
  not NOT_1947(g4493,I8543);
  not NOT_1948(g7764,I14163);
  not NOT_1949(g6351,I11380);
  not NOT_1950(g6648,I11926);
  not NOT_1951(g6875,I12496);
  not NOT_1952(g7546,I13822);
  not NOT_1953(g3865,g2944);
  not NOT_1954(I10384,g5193);
  not NOT_1955(g6655,I11945);
  not NOT_1956(g5445,g5059);
  not NOT_1957(g5173,I9645);
  not NOT_1958(I11317,g5787);
  not NOT_1959(g3604,g2407);
  not NOT_1960(I13317,g7211);
  not NOT_1961(g5491,g4918);
  not NOT_1962(g3498,g1616);
  not NOT_1963(I14067,g7550);
  not NOT_1964(I14094,g7593);
  not NOT_1965(g4381,g3466);
  not NOT_1966(g8649,I14743);
  not NOT_1967(g6010,I10608);
  not NOT_1968(g3833,I7302);
  not NOT_1969(I11129,g5418);
  not NOT_1970(g2872,I6590);
  not NOT_1971(g1924,g174);
  not NOT_1972(g5169,I9633);
  not NOT_1973(g4685,I8952);
  not NOT_1974(g4197,g3591);
  not NOT_1975(I10801,g5463);
  not NOT_1976(g6410,I11533);
  not NOT_1977(g7224,I13164);
  not NOT_1978(I7520,g2734);
  not NOT_1979(g4021,g3131);
  not NOT_1980(g5007,I9336);
  not NOT_1981(I13057,g6968);
  not NOT_1982(I14801,g8608);
  not NOT_1983(g2652,I6440);
  not NOT_1984(g1779,g612);
  not NOT_1985(g2057,I5868);
  not NOT_1986(I7640,g3062);
  not NOT_1987(I12124,g5847);
  not NOT_1988(I12678,g6516);
  not NOT_1989(g6884,I12523);
  not NOT_1990(g2843,I6571);
  not NOT_1991(g7120,I12948);
  not NOT_1992(g5059,I9419);
  not NOT_1993(g6839,I12388);
  not NOT_1994(g2457,g24);
  not NOT_1995(g5578,g4841);
  not NOT_1996(g5868,I10555);
  not NOT_1997(g7320,I13388);
  not NOT_1998(g2989,g1843);
  not NOT_1999(g3539,g2424);
  not NOT_2000(g3896,I7473);
  not NOT_2001(I11245,g6143);
  not NOT_2002(g5459,g4882);
  not NOT_2003(I14019,g7480);
  not NOT_2004(g2393,I6267);
  not NOT_2005(g5718,g4841);
  not NOT_2006(I12460,g6674);
  not NOT_2007(I12939,g7022);
  not NOT_2008(I11323,g5808);
  not NOT_2009(g1977,g1357);
  not NOT_2010(I11299,g5786);
  not NOT_2011(I13323,g7145);
  not NOT_2012(I14196,g7534);
  not NOT_2013(I13299,g7163);
  not NOT_2014(I14695,g8016);
  not NOT_2015(g7277,I13267);
  not NOT_2016(g1588,g741);
  not NOT_2017(I11533,g5847);
  not NOT_2018(g2834,I6564);
  not NOT_2019(g2971,I6723);
  not NOT_2020(I13533,g7220);
  not NOT_2021(g8063,I14334);
  not NOT_2022(g5582,g4969);
  not NOT_2023(I15405,g8902);
  not NOT_2024(g6278,I11129);
  not NOT_2025(g8463,g8094);
  not NOT_2026(g2686,g1667);
  not NOT_2027(g6372,I11443);
  not NOT_2028(g7789,I14224);
  not NOT_2029(g5261,g4748);
  not NOT_2030(g3019,g2007);
  not NOT_2031(g9132,I15770);
  not NOT_2032(g5793,I10418);
  not NOT_2033(I12065,g5897);
  not NOT_2034(I8202,g3560);
  not NOT_2035(g9332,g9322);
  not NOT_2036(g6618,g6003);
  not NOT_2037(g1665,g1467);
  not NOT_2038(g6143,I10796);
  not NOT_2039(g7516,I13728);
  not NOT_2040(I7765,g2595);
  not NOT_2041(g6343,I11356);
  not NOT_2042(g4562,g3466);
  not NOT_2043(g6235,I11034);
  not NOT_2044(g5015,I9347);
  not NOT_2045(g3052,g2096);
  not NOT_2046(g9209,g9199);
  not NOT_2047(g9353,I16107);
  not NOT_2048(I7911,g2767);
  not NOT_2049(I10457,g5218);
  not NOT_2050(I8094,g2976);
  not NOT_2051(g7771,I14184);
  not NOT_2052(I14457,g8093);
  not NOT_2053(g6566,I11740);
  not NOT_2054(g4631,I8808);
  not NOT_2055(I13737,g7446);
  not NOT_2056(g372,I5359);
  not NOT_2057(I15583,g8986);
  not NOT_2058(g7299,I13329);
  not NOT_2059(g4257,I8190);
  not NOT_2060(g6693,I12011);
  not NOT_2061(g6134,g5428);
  not NOT_2062(g8619,I14695);
  not NOT_2063(g7547,I13825);
  not NOT_2064(g6334,I11329);
  not NOT_2065(g4301,I8264);
  not NOT_2066(g5246,I9760);
  not NOT_2067(g2625,g1570);
  not NOT_2068(g8872,I15202);
  not NOT_2069(g2232,I5957);
  not NOT_2070(g4605,I8730);
  not NOT_2071(g3086,g1852);
  not NOT_2072(g2253,g1323);
  not NOT_2073(g2938,g2347);
  not NOT_2074(g3728,g2202);
  not NOT_2075(I14001,g7433);
  not NOT_2076(I13261,g7041);
  not NOT_2077(I11880,g5748);
  not NOT_2078(g6555,I11729);
  not NOT_2079(g6804,I12283);
  not NOT_2080(I7473,g3546);
  not NOT_2081(g2909,g2291);
  not NOT_2082(I6946,g1887);
  not NOT_2083(I10256,g5401);
  not NOT_2084(g6792,I12247);
  not NOT_2085(I11512,g5874);
  not NOT_2086(g1732,g1439);
  not NOT_2087(I9675,g4807);
  not NOT_2088(I13512,g7138);
  not NOT_2089(g3881,g2969);
  not NOT_2090(I5383,g647);
  not NOT_2091(I10280,g5488);
  not NOT_2092(g8971,I15417);
  not NOT_2093(g7738,I14085);
  not NOT_2094(g4585,g2925);
  not NOT_2095(I8264,g3653);
  not NOT_2096(g6621,I11855);
  not NOT_2097(g1944,I5817);
  not NOT_2098(g3897,g3131);
  not NOT_2099(g4041,g2605);
  not NOT_2100(I12915,g7000);
  not NOT_2101(g9092,I15666);
  not NOT_2102(I8360,g1186);
  not NOT_2103(g6313,I11266);
  not NOT_2104(g7078,g6683);
  not NOT_2105(g7340,I13438);
  not NOT_2106(I7377,g3189);
  not NOT_2107(I10157,g5109);
  not NOT_2108(I13831,g7322);
  not NOT_2109(I6036,g130);
  not NOT_2110(I14157,g7547);
  not NOT_2111(I12277,g6681);
  not NOT_2112(I6178,g1220);
  not NOT_2113(g4673,I8928);
  not NOT_2114(g6202,I10949);
  not NOT_2115(g8670,I14804);
  not NOT_2116(I9684,g4813);
  not NOT_2117(g7035,g6543);
  not NOT_2118(I13499,g7134);
  not NOT_2119(I15803,g9148);
  not NOT_2120(I9639,g4685);
  not NOT_2121(g7517,I13731);
  not NOT_2122(I7287,g2561);
  not NOT_2123(g6094,I10716);
  not NOT_2124(I14231,g7566);
  not NOT_2125(I9791,g4779);
  not NOT_2126(I6831,g2185);
  not NOT_2127(g5028,I9372);
  not NOT_2128(g4669,I8922);
  not NOT_2129(g1565,g649);
  not NOT_2130(I8724,g3927);
  not NOT_2131(g5671,I10160);
  not NOT_2132(I11722,g5772);
  not NOT_2133(I12782,g6463);
  not NOT_2134(I13722,g7442);
  not NOT_2135(I16090,g9336);
  not NOT_2136(I6805,g1603);
  not NOT_2137(g3635,g1949);
  not NOT_2138(I13924,g7365);
  not NOT_2139(I5633,g891);
  not NOT_2140(g1681,g929);
  not NOT_2141(g6776,I12199);
  not NOT_2142(I7781,g2605);
  not NOT_2143(I6422,g1805);
  not NOT_2144(g6593,I11793);
  not NOT_2145(g4890,g4075);
  not NOT_2146(I12352,g6752);
  not NOT_2147(I13432,g7280);
  not NOT_2148(g2525,I6354);
  not NOT_2149(g3801,I7262);
  not NOT_2150(I14763,g7834);
  not NOT_2151(I13271,g7067);
  not NOT_2152(g2645,I6419);
  not NOT_2153(I8835,g3954);
  not NOT_2154(g5826,I10503);
  not NOT_2155(I12418,g6572);
  not NOT_2156(I7797,g3019);
  not NOT_2157(g8606,I14683);
  not NOT_2158(I12170,g5956);
  not NOT_2159(g4011,I7762);
  not NOT_2160(I11461,g6094);
  not NOT_2161(g9076,I15622);
  not NOT_2162(g5741,I10280);
  not NOT_2163(g7110,I12918);
  not NOT_2164(I5732,g859);
  not NOT_2165(g6264,g5403);
  not NOT_2166(g7310,I13362);
  not NOT_2167(I11031,g5335);
  not NOT_2168(I13031,g6984);
  not NOT_2169(g5638,g4748);
  not NOT_2170(g6360,I11407);
  not NOT_2171(g2879,I6597);
  not NOT_2172(I13199,g7025);
  not NOT_2173(I11736,g6076);
  not NOT_2174(I11887,g5918);
  not NOT_2175(g9375,I16151);
  not NOT_2176(I7344,g2964);
  not NOT_2177(g2962,g2382);
  not NOT_2178(g5609,g4748);
  not NOT_2179(I15003,g8633);
  not NOT_2180(I8799,g3951);
  not NOT_2181(g2659,g1655);
  not NOT_2182(g6050,g5246);
  not NOT_2183(I12167,g5939);
  not NOT_2184(g2506,I6341);
  not NOT_2185(g1820,g621);
  not NOT_2186(I6437,g1784);
  not NOT_2187(I11696,g5971);
  not NOT_2188(g7236,g6944);
  not NOT_2189(I6302,g1313);
  not NOT_2190(g3091,g1603);
  not NOT_2191(I13843,g7326);
  not NOT_2192(I16026,g9267);
  not NOT_2193(g7762,I14157);
  not NOT_2194(g3491,g1800);
  not NOT_2195(g4080,I7867);
  not NOT_2196(I14076,g7577);
  not NOT_2197(I14085,g7583);
  not NOT_2198(g4573,g2911);
  not NOT_2199(I11764,g6056);
  not NOT_2200(g5758,I10347);
  not NOT_2201(I13764,g7479);
  not NOT_2202(g6724,I12088);
  not NOT_2203(I11365,g5826);
  not NOT_2204(g2275,g990);
  not NOT_2205(g2311,I6090);
  not NOT_2206(I9539,g4018);
  not NOT_2207(g6179,I10896);
  not NOT_2208(I13365,g7267);
  not NOT_2209(g5466,g4890);
  not NOT_2210(g4713,I9014);
  not NOT_2211(I10243,g5026);
  not NOT_2212(g6379,I11464);
  not NOT_2213(I11132,g5624);
  not NOT_2214(g7590,I13915);
  not NOT_2215(g9184,I15830);
  not NOT_2216(I13869,g7338);
  not NOT_2217(I5565,g1296);
  not NOT_2218(g2615,g1563);
  not NOT_2219(g6878,I12505);
  not NOT_2220(g5165,I9621);
  not NOT_2221(g4569,g2906);
  not NOT_2222(g5571,I10032);
  not NOT_2223(g3920,g3097);
  not NOT_2224(I12022,g5874);
  not NOT_2225(g3578,I7053);
  not NOT_2226(g3868,g2948);
  not NOT_2227(g2174,g1319);
  not NOT_2228(g6289,I11194);
  not NOT_2229(g6777,I12202);
  not NOT_2230(I8802,g3963);
  not NOT_2231(g6658,g6224);
  not NOT_2232(g2374,I6220);
  not NOT_2233(g5448,g5137);
  not NOT_2234(g1922,g1251);
  not NOT_2235(I9162,g4272);
  not NOT_2236(g7556,I13846);
  not NOT_2237(I13161,g7080);
  not NOT_2238(I10773,g5708);
  not NOT_2239(g5055,g4477);
  not NOT_2240(I12313,g6730);
  not NOT_2241(g6835,I12376);
  not NOT_2242(g2985,I6733);
  not NOT_2243(I9419,g3916);
  not NOT_2244(I10268,g5471);
  not NOT_2245(g1581,g710);
  not NOT_2246(g5827,I10506);
  not NOT_2247(I12748,g6585);
  not NOT_2248(g6882,I12517);
  not NOT_2249(I6042,g237);
  not NOT_2250(I15651,g9056);
  not NOT_2251(I15672,g9047);
  not NOT_2252(g3582,g2407);
  not NOT_2253(g2284,I6036);
  not NOT_2254(I5914,g1097);
  not NOT_2255(I13225,g7095);
  not NOT_2256(g7064,I12829);
  not NOT_2257(g2239,I5978);
  not NOT_2258(I7314,g2916);
  not NOT_2259(I10180,g4721);
  not NOT_2260(I16148,g9368);
  not NOT_2261(g1597,g973);
  not NOT_2262(g9077,I15625);
  not NOT_2263(g2180,g1318);
  not NOT_2264(g5846,g5367);
  not NOT_2265(g2380,I6242);
  not NOT_2266(I13258,g6907);
  not NOT_2267(I12900,g6947);
  not NOT_2268(I7870,g2827);
  not NOT_2269(I8901,g4122);
  not NOT_2270(g2832,g2184);
endmodule