// Verilog
// c3540
// Ninputs 50
// Noutputs 22
// NtotalGates 1669
// BUFF1 223
// NOT1 490
// OR2 35
// AND2 410
// NAND2 274
// NAND3 17
// AND3 76
// NOR2 25
// AND4 10
// NAND4 7
// OR3 56
// NOR3 27
// AND5 2
// NOR8 16
// OR4 1

module c3540 (N1,N13,N20,N33,N41,N45,N50,N58,N68,N77,
              N87,N97,N107,N116,N124,N125,N128,N132,N137,N143,
              N150,N159,N169,N179,N190,N200,N213,N222,N223,N226,
              N232,N238,N244,N250,N257,N264,N270,N274,N283,N294,
              N303,N311,N317,N322,N326,N329,N330,N343,N349,N350,
              N1713,N1947,N3195,N3833,N3987,N4028,N4145,N4589,N4667,N4815,
              N4944,N5002,N5045,N5047,N5078,N5102,N5120,N5121,N5192,N5231,
              N5360,N5361,clk);

input N1,N13,N20,N33,N41,N45,N50,N58,N68,N77,
      N87,N97,N107,N116,N124,N125,N128,N132,N137,N143,
      N150,N159,N169,N179,N190,N200,N213,N222,N223,N226,
      N232,N238,N244,N250,N257,N264,N270,N274,N283,N294,
      N303,N311,N317,N322,N326,N329,N330,N343,N349,N350,clk;

output N1713,N1947,N3195,N3833,N3987,N4028,N4145,N4589,N4667,N4815,
       N4944,N5002,N5045,N5047,N5078,N5102,N5120,N5121,N5192,N5231,
       N5360,N5361;

wire N655,N665,N670,N679,N683,N686,N690,N699,N702,N706,
     N715,N724,N727,N736,N740,N749,N753,N763,N768,N769,
     N772,N779,N782,N786,N793,N794,N798,N803,N820,N821,
     N825,N829,N832,N835,N836,N839,N842,N845,N848,N851,
     N854,N858,N861,N864,N867,N870,N874,N877,N880,N883,
     N886,N889,N890,N891,N892,N895,N896,N913,N914,N915,
     N916,N917,N920,N923,N926,N929,N932,N935,N938,N941,
     N944,N947,N950,N953,N956,N959,N962,N965,N1067,N1117,
     N1179,N1196,N1197,N1202,N1219,N1250,N1251,N1252,N1253,N1254,
     N1255,N1256,N1257,N1258,N1259,N1260,N1261,N1262,N1263,N1264,
     N1267,N1268,N1271,N1272,N1273,N1276,N1279,N1298,N1302,N1306,
     N1315,N1322,N1325,N1328,N1331,N1334,N1337,N1338,N1339,N1340,
     N1343,N1344,N1345,N1346,N1347,N1348,N1349,N1350,N1351,N1352,
     N1353,N1358,N1363,N1366,N1369,N1384,N1401,N1402,N1403,N1404,
     N1405,N1406,N1407,N1408,N1409,N1426,N1427,N1452,N1459,N1460,
     N1461,N1464,N1467,N1468,N1469,N1470,N1471,N1474,N1475,N1478,
     N1481,N1484,N1487,N1490,N1493,N1496,N1499,N1502,N1505,N1507,
     N1508,N1509,N1510,N1511,N1512,N1520,N1562,N1579,N1580,N1581,
     N1582,N1583,N1584,N1585,N1586,N1587,N1588,N1589,N1590,N1591,
     N1592,N1593,N1594,N1595,N1596,N1597,N1598,N1599,N1600,N1643,
     N1644,N1645,N1646,N1647,N1648,N1649,N1650,N1667,N1670,N1673,
     N1674,N1675,N1676,N1677,N1678,N1679,N1680,N1691,N1692,N1693,
     N1694,N1714,N1715,N1718,N1721,N1722,N1725,N1726,N1727,N1728,
     N1729,N1730,N1731,N1735,N1736,N1737,N1738,N1747,N1756,N1761,
     N1764,N1765,N1766,N1767,N1768,N1769,N1770,N1787,N1788,N1789,
     N1790,N1791,N1792,N1793,N1794,N1795,N1796,N1797,N1798,N1799,
     N1800,N1801,N1802,N1803,N1806,N1809,N1812,N1815,N1818,N1821,
     N1824,N1833,N1842,N1843,N1844,N1845,N1846,N1847,N1848,N1849,
     N1850,N1851,N1852,N1853,N1854,N1855,N1856,N1857,N1858,N1859,
     N1860,N1861,N1862,N1863,N1864,N1869,N1870,N1873,N1874,N1875,
     N1878,N1879,N1880,N1883,N1884,N1885,N1888,N1889,N1890,N1893,
     N1894,N1895,N1898,N1899,N1900,N1903,N1904,N1905,N1908,N1909,
     N1912,N1913,N1917,N1922,N1926,N1930,N1933,N1936,N1939,N1940,
     N1941,N1942,N1943,N1944,N1945,N1946,N1960,N1961,N1966,N1981,
     N1982,N1983,N1986,N1987,N1988,N1989,N1990,N1991,N2022,N2023,
     N2024,N2025,N2026,N2027,N2028,N2029,N2030,N2031,N2032,N2033,
     N2034,N2035,N2036,N2037,N2038,N2043,N2052,N2057,N2068,N2073,
     N2078,N2083,N2088,N2093,N2098,N2103,N2121,N2122,N2123,N2124,
     N2125,N2126,N2127,N2128,N2133,N2134,N2135,N2136,N2137,N2138,
     N2139,N2141,N2142,N2143,N2144,N2145,N2146,N2147,N2148,N2149,
     N2150,N2151,N2152,N2153,N2154,N2155,N2156,N2157,N2158,N2175,
     N2178,N2179,N2180,N2181,N2183,N2184,N2185,N2188,N2191,N2194,
     N2197,N2200,N2203,N2206,N2209,N2210,N2211,N2212,N2221,N2230,
     N2231,N2232,N2233,N2234,N2235,N2236,N2237,N2238,N2239,N2240,
     N2241,N2242,N2243,N2244,N2245,N2270,N2277,N2282,N2287,N2294,
     N2299,N2304,N2307,N2310,N2313,N2316,N2319,N2322,N2325,N2328,
     N2331,N2334,N2341,N2342,N2347,N2348,N2349,N2350,N2351,N2352,
     N2353,N2354,N2355,N2374,N2375,N2376,N2379,N2398,N2417,N2418,
     N2419,N2420,N2421,N2422,N2425,N2426,N2427,N2430,N2431,N2432,
     N2435,N2436,N2437,N2438,N2439,N2440,N2443,N2444,N2445,N2448,
     N2449,N2450,N2467,N2468,N2469,N2470,N2471,N2474,N2475,N2476,
     N2477,N2478,N2481,N2482,N2483,N2486,N2487,N2488,N2497,N2506,
     N2515,N2524,N2533,N2542,N2551,N2560,N2569,N2578,N2587,N2596,
     N2605,N2614,N2623,N2632,N2633,N2634,N2635,N2636,N2637,N2638,
     N2639,N2640,N2641,N2642,N2643,N2644,N2645,N2646,N2647,N2648,
     N2652,N2656,N2659,N2662,N2666,N2670,N2673,N2677,N2681,N2684,
     N2688,N2692,N2697,N2702,N2706,N2710,N2715,N2719,N2723,N2728,
     N2729,N2730,N2731,N2732,N2733,N2734,N2735,N2736,N2737,N2738,
     N2739,N2740,N2741,N2742,N2743,N2744,N2745,N2746,N2748,N2749,
     N2750,N2751,N2754,N2755,N2756,N2757,N2758,N2761,N2764,N2768,
     N2769,N2898,N2899,N2900,N2901,N2962,N2966,N2967,N2970,N2973,
     N2977,N2980,N2984,N2985,N2986,N2987,N2988,N2989,N2990,N2991,
     N2992,N2993,N2994,N2995,N2996,N2997,N2998,N2999,N3000,N3001,
     N3002,N3003,N3004,N3005,N3006,N3007,N3008,N3009,N3010,N3011,
     N3012,N3013,N3014,N3015,N3016,N3017,N3018,N3019,N3020,N3021,
     N3022,N3023,N3024,N3025,N3026,N3027,N3028,N3029,N3030,N3031,
     N3032,N3033,N3034,N3035,N3036,N3037,N3038,N3039,N3040,N3041,
     N3042,N3043,N3044,N3045,N3046,N3047,N3048,N3049,N3050,N3051,
     N3052,N3053,N3054,N3055,N3056,N3057,N3058,N3059,N3060,N3061,
     N3062,N3063,N3064,N3065,N3066,N3067,N3068,N3069,N3070,N3071,
     N3072,N3073,N3074,N3075,N3076,N3077,N3078,N3079,N3080,N3081,
     N3082,N3083,N3084,N3085,N3086,N3087,N3088,N3089,N3090,N3091,
     N3092,N3093,N3094,N3095,N3096,N3097,N3098,N3099,N3100,N3101,
     N3102,N3103,N3104,N3105,N3106,N3107,N3108,N3109,N3110,N3111,
     N3112,N3115,N3118,N3119,N3122,N3125,N3128,N3131,N3134,N3135,
     N3138,N3141,N3142,N3145,N3148,N3149,N3152,N3155,N3158,N3161,
     N3164,N3165,N3168,N3171,N3172,N3175,N3178,N3181,N3184,N3187,
     N3190,N3191,N3192,N3193,N3194,N3196,N3206,N3207,N3208,N3209,
     N3210,N3211,N3212,N3213,N3214,N3215,N3216,N3217,N3218,N3219,
     N3220,N3221,N3222,N3223,N3224,N3225,N3226,N3227,N3228,N3229,
     N3230,N3231,N3232,N3233,N3234,N3235,N3236,N3237,N3238,N3239,
     N3240,N3241,N3242,N3243,N3244,N3245,N3246,N3247,N3248,N3249,
     N3250,N3251,N3252,N3253,N3254,N3255,N3256,N3257,N3258,N3259,
     N3260,N3261,N3262,N3263,N3264,N3265,N3266,N3267,N3268,N3269,
     N3270,N3271,N3272,N3273,N3274,N3275,N3276,N3277,N3278,N3279,
     N3280,N3281,N3282,N3283,N3284,N3285,N3286,N3287,N3288,N3289,
     N3290,N3291,N3292,N3293,N3294,N3295,N3296,N3297,N3298,N3299,
     N3300,N3301,N3302,N3303,N3304,N3305,N3306,N3307,N3308,N3309,
     N3310,N3311,N3312,N3313,N3314,N3315,N3316,N3317,N3318,N3319,
     N3320,N3321,N3322,N3323,N3324,N3325,N3326,N3327,N3328,N3329,
     N3330,N3331,N3332,N3333,N3334,N3383,N3384,N3387,N3388,N3389,
     N3390,N3391,N3392,N3393,N3394,N3395,N3396,N3397,N3398,N3399,
     N3400,N3401,N3402,N3403,N3404,N3405,N3406,N3407,N3410,N3413,
     N3414,N3415,N3419,N3423,N3426,N3429,N3430,N3431,N3434,N3437,
     N3438,N3439,N3442,N3445,N3446,N3447,N3451,N3455,N3458,N3461,
     N3462,N3463,N3466,N3469,N3470,N3471,N3472,N3475,N3478,N3481,
     N3484,N3487,N3490,N3493,N3496,N3499,N3502,N3505,N3508,N3511,
     N3514,N3517,N3520,N3523,N3534,N3535,N3536,N3537,N3538,N3539,
     N3540,N3541,N3542,N3543,N3544,N3545,N3546,N3547,N3548,N3549,
     N3550,N3551,N3552,N3557,N3568,N3573,N3578,N3589,N3594,N3605,
     N3626,N3627,N3628,N3629,N3630,N3631,N3632,N3633,N3634,N3635,
     N3636,N3637,N3638,N3639,N3640,N3641,N3642,N3643,N3644,N3645,
     N3648,N3651,N3652,N3653,N3654,N3657,N3658,N3661,N3662,N3663,
     N3664,N3667,N3670,N3671,N3672,N3673,N3676,N3677,N3680,N3681,
     N3682,N3685,N3686,N3687,N3688,N3689,N3690,N3693,N3694,N3695,
     N3696,N3697,N3700,N3703,N3704,N3705,N3706,N3707,N3708,N3711,
     N3712,N3713,N3714,N3715,N3716,N3717,N3718,N3719,N3720,N3721,
     N3731,N3734,N3740,N3743,N3753,N3756,N3762,N3765,N3766,N3773,
     N3774,N3775,N3776,N3777,N3778,N3779,N3780,N3786,N3789,N3800,
     N3803,N3809,N3812,N3815,N3818,N3821,N3824,N3827,N3830,N3834,
     N3835,N3838,N3845,N3850,N3855,N3858,N3861,N3865,N3868,N3884,
     N3885,N3894,N3895,N3898,N3899,N3906,N3911,N3912,N3913,N3916,
     N3917,N3920,N3921,N3924,N3925,N3926,N3930,N3931,N3932,N3935,
     N3936,N3937,N3940,N3947,N3948,N3950,N3953,N3956,N3959,N3962,
     N3965,N3968,N3971,N3974,N3977,N3980,N3983,N3992,N3996,N4013,
     N4029,N4030,N4031,N4032,N4033,N4034,N4035,N4042,N4043,N4044,
     N4045,N4046,N4047,N4048,N4049,N4050,N4051,N4052,N4053,N4054,
     N4055,N4056,N4057,N4058,N4059,N4062,N4065,N4066,N4067,N4070,
     N4073,N4074,N4075,N4076,N4077,N4078,N4079,N4080,N4085,N4086,
     N4088,N4090,N4091,N4094,N4098,N4101,N4104,N4105,N4106,N4107,
     N4108,N4109,N4110,N4111,N4112,N4113,N4114,N4115,N4116,N4119,
     N4122,N4123,N4126,N4127,N4128,N4139,N4142,N4146,N4147,N4148,
     N4149,N4150,N4151,N4152,N4153,N4154,N4161,N4167,N4174,N4182,
     N4186,N4189,N4190,N4191,N4192,N4193,N4194,N4195,N4196,N4197,
     N4200,N4203,N4209,N4213,N4218,N4223,N4238,N4239,N4241,N4242,
     N4247,N4251,N4252,N4253,N4254,N4255,N4256,N4257,N4258,N4283,
     N4284,N4287,N4291,N4295,N4296,N4299,N4303,N4304,N4305,N4310,
     N4316,N4317,N4318,N4319,N4322,N4325,N4326,N4327,N4328,N4329,
     N4330,N4331,N4335,N4338,N4341,N4344,N4347,N4350,N4353,N4356,
     N4359,N4362,N4365,N4368,N4371,N4376,N4377,N4387,N4390,N4393,
     N4398,N4413,N4416,N4421,N4427,N4430,N4435,N4442,N4443,N4446,
     N4447,N4448,N4452,N4458,N4461,N4462,N4463,N4464,N4465,N4468,
     N4472,N4475,N4479,N4484,N4486,N4487,N4491,N4493,N4496,N4497,
     N4498,N4503,N4506,N4507,N4508,N4509,N4510,N4511,N4515,N4526,
     N4527,N4528,N4529,N4530,N4531,N4534,N4537,N4540,N4545,N4549,
     N4552,N4555,N4558,N4559,N4562,N4563,N4564,N4568,N4569,N4572,
     N4573,N4576,N4581,N4584,N4587,N4588,N4593,N4596,N4597,N4599,
     N4602,N4603,N4608,N4613,N4616,N4619,N4623,N4628,N4629,N4630,
     N4635,N4636,N4640,N4641,N4642,N4643,N4644,N4647,N4650,N4656,
     N4659,N4664,N4668,N4669,N4670,N4673,N4674,N4675,N4676,N4677,
     N4678,N4679,N4687,N4688,N4691,N4694,N4697,N4700,N4704,N4705,
     N4706,N4707,N4708,N4711,N4716,N4717,N4721,N4722,N4726,N4727,
     N4730,N4733,N4740,N4743,N4747,N4748,N4749,N4750,N4753,N4754,
     N4755,N4756,N4757,N4769,N4772,N4775,N4778,N4786,N4787,N4788,
     N4789,N4794,N4797,N4800,N4805,N4808,N4812,N4816,N4817,N4818,
     N4822,N4823,N4826,N4829,N4830,N4831,N4838,N4844,N4847,N4850,
     N4854,N4859,N4860,N4868,N4870,N4872,N4873,N4876,N4880,N4885,
     N4889,N4895,N4896,N4897,N4898,N4899,N4900,N4901,N4902,N4904,
     N4905,N4906,N4907,N4913,N4916,N4920,N4921,N4924,N4925,N4926,
     N4928,N4929,N4930,N4931,N4937,N4940,N4946,N4949,N4950,N4951,
     N4952,N4953,N4954,N4957,N4964,N4965,N4968,N4969,N4970,N4973,
     N4978,N4979,N4980,N4981,N4982,N4983,N4984,N4985,N4988,N4991,
     N4996,N4999,N5007,N5010,N5013,N5018,N5021,N5026,N5029,N5030,
     N5039,N5042,N5046,N5050,N5055,N5058,N5061,N5066,N5070,N5080,
     N5085,N5094,N5095,N5097,N5103,N5108,N5109,N5110,N5111,N5114,
     N5117,N5122,N5125,N5128,N5133,N5136,N5139,N5145,N5151,N5154,
     N5159,N5160,N5163,N5166,N5173,N5174,N5177,N5182,N5183,N5184,
     N5188,N5193,N5196,N5197,N5198,N5199,N5201,N5203,N5205,N5209,
     N5212,N5215,N5217,N5219,N5220,N5221,N5222,N5223,N5224,N5225,
     N5228,N5232,N5233,N5234,N5235,N5236,N5240,N5242,N5243,N5245,
     N5246,N5250,N5253,N5254,N5257,N5258,N5261,N5266,N5269,N5277,
     N5278,N5279,N5283,N5284,N5285,N5286,N5289,N5292,N5295,N5298,
     N5303,N5306,N5309,N5312,N5313,N5322,N5323,N5324,N5327,N5332,
     N5335,N5340,N5341,N5344,N5345,N5348,N5349,N5350,N5351,N5352,
     N5353,N5354,N5355,N5356,N5357,N5358,N5359;

buf BUFF1_1 (N655, N50);
not NOT1_2 (N665, N50);
buf BUFF1_3 (N670, N58);
not NOT1_4 (N679, N58);
buf BUFF1_5 (N683, N68);
not NOT1_6 (N686, N68);
buf BUFF1_7 (N690, N68);
buf BUFF1_8 (N699, N77);
not NOT1_9 (N702, N77);
buf BUFF1_10 (N706, N77);
buf BUFF1_11 (N715, N87);
not NOT1_12 (N724, N87);
buf BUFF1_13 (N727, N97);
not NOT1_14 (N736, N97);
buf BUFF1_15 (N740, N107);
not NOT1_16 (N749, N107);
buf BUFF1_17 (N753, N116);
not NOT1_18 (N763, N116);
or OR2_19 (N768, N257, N264);
not NOT1_20 (N769, N1);
buf BUFF1_21 (N772, N1);
not NOT1_22 (N779, N1);
buf BUFF1_23 (N782, N13);
not NOT1_24 (N786, N13);
and AND2_25 (N793, N13, N20);
not NOT1_26 (N794, N20);
buf BUFF1_27 (N798, N20);
not NOT1_28 (N803, N20);
not NOT1_29 (N820, N33);
buf BUFF1_30 (N821, N33);
not NOT1_31 (N825, N33);
and AND2_32 (N829, N33, N41);
not NOT1_33 (N832, N41);
or OR2_34 (N835, N41, N45);
buf BUFF1_35 (N836, N45);
not NOT1_36 (N839, N45);
not NOT1_37 (N842, N50);
buf BUFF1_38 (N845, N58);
not NOT1_39 (N848, N58);
buf BUFF1_40 (N851, N68);
not NOT1_41 (N854, N68);
buf BUFF1_42 (N858, N87);
not NOT1_43 (N861, N87);
buf BUFF1_44 (N864, N97);
not NOT1_45 (N867, N97);
not NOT1_46 (N870, N107);
buf BUFF1_47 (N874, N1);
buf BUFF1_48 (N877, N68);
buf BUFF1_49 (N880, N107);
not NOT1_50 (N883, N20);
buf BUFF1_51 (N886, N190);
not NOT1_52 (N889, N200);
and AND2_53 (N890, N20, N200);
nand NAND2_54 (N891, N20, N200);
and AND2_55 (N892, N20, N179);
not NOT1_56 (N895, N20);
or OR2_57 (N896, N349, N33);
nand NAND2_58 (N913, N1, N13);
nand NAND3_59 (N914, N1, N20, N33);
not NOT1_60 (N915, N20);
not NOT1_61 (N916, N33);
buf BUFF1_62 (N917, N179);
not NOT1_63 (N920, N213);
buf BUFF1_64 (N923, N343);
buf BUFF1_65 (N926, N226);
buf BUFF1_66 (N929, N232);
buf BUFF1_67 (N932, N238);
buf BUFF1_68 (N935, N244);
buf BUFF1_69 (N938, N250);
buf BUFF1_70 (N941, N257);
buf BUFF1_71 (N944, N264);
buf BUFF1_72 (N947, N270);
buf BUFF1_73 (N950, N50);
buf BUFF1_74 (N953, N58);
buf BUFF1_75 (N956, N58);
buf BUFF1_76 (N959, N97);
buf BUFF1_77 (N962, N97);
buf BUFF1_78 (N965, N330);
and AND2_79 (N1067, N250, N768);
or OR2_80 (N1117, N820, N20);
or OR2_81 (N1179, N895, N169);
not NOT1_82 (N1196, N793);
or OR2_83 (N1197, N915, N1);
and AND2_84 (N1202, N913, N914);
or OR2_85 (N1219, N916, N1);
and AND3_86 (N1250, N842, N848, N854);
nand NAND2_87 (N1251, N226, N655);
nand NAND2_88 (N1252, N232, N670);
nand NAND2_89 (N1253, N238, N690);
nand NAND2_90 (N1254, N244, N706);
nand NAND2_91 (N1255, N250, N715);
nand NAND2_92 (N1256, N257, N727);
nand NAND2_93 (N1257, N264, N740);
nand NAND2_94 (N1258, N270, N753);
not NOT1_95 (N1259, N926);
not NOT1_96 (N1260, N929);
not NOT1_97 (N1261, N932);
not NOT1_98 (N1262, N935);
nand NAND2_99 (N1263, N679, N686);
nand NAND2_100 (N1264, N736, N749);
nand NAND2_101 (N1267, N683, N699);
buf BUFF1_102 (N1268, N665);
not NOT1_103 (N1271, N953);
not NOT1_104 (N1272, N959);
buf BUFF1_105 (N1273, N839);
buf BUFF1_106 (N1276, N839);
buf BUFF1_107 (N1279, N782);
buf BUFF1_108 (N1298, N825);
buf BUFF1_109 (N1302, N832);
and AND2_110 (N1306, N779, N835);
and AND3_111 (N1315, N779, N836, N832);
and AND2_112 (N1322, N769, N836);
and AND3_113 (N1325, N772, N786, N798);
nand NAND3_114 (N1328, N772, N786, N798);
nand NAND2_115 (N1331, N772, N786);
buf BUFF1_116 (N1334, N874);
nand NAND3_117 (N1337, N782, N794, N45);
nand NAND3_118 (N1338, N842, N848, N854);
not NOT1_119 (N1339, N956);
and AND3_120 (N1340, N861, N867, N870);
nand NAND3_121 (N1343, N861, N867, N870);
not NOT1_122 (N1344, N962);
not NOT1_123 (N1345, N803);
not NOT1_124 (N1346, N803);
not NOT1_125 (N1347, N803);
not NOT1_126 (N1348, N803);
not NOT1_127 (N1349, N803);
not NOT1_128 (N1350, N803);
not NOT1_129 (N1351, N803);
not NOT1_130 (N1352, N803);
or OR2_131 (N1353, N883, N886);
nor NOR2_132 (N1358, N883, N886);
buf BUFF1_133 (N1363, N892);
not NOT1_134 (N1366, N892);
buf BUFF1_135 (N1369, N821);
buf BUFF1_136 (N1384, N825);
not NOT1_137 (N1401, N896);
not NOT1_138 (N1402, N896);
not NOT1_139 (N1403, N896);
not NOT1_140 (N1404, N896);
not NOT1_141 (N1405, N896);
not NOT1_142 (N1406, N896);
not NOT1_143 (N1407, N896);
not NOT1_144 (N1408, N896);
or OR2_145 (N1409, N1, N1196);
not NOT1_146 (N1426, N829);
not NOT1_147 (N1427, N829);
and AND3_148 (N1452, N769, N782, N794);
not NOT1_149 (N1459, N917);
not NOT1_150 (N1460, N965);
or OR2_151 (N1461, N920, N923);
nor NOR2_152 (N1464, N920, N923);
not NOT1_153 (N1467, N938);
not NOT1_154 (N1468, N941);
not NOT1_155 (N1469, N944);
not NOT1_156 (N1470, N947);
buf BUFF1_157 (N1471, N679);
not NOT1_158 (N1474, N950);
buf BUFF1_159 (N1475, N686);
buf BUFF1_160 (N1478, N702);
buf BUFF1_161 (N1481, N724);
buf BUFF1_162 (N1484, N736);
buf BUFF1_163 (N1487, N749);
buf BUFF1_164 (N1490, N763);
buf BUFF1_165 (N1493, N877);
buf BUFF1_166 (N1496, N877);
buf BUFF1_167 (N1499, N880);
buf BUFF1_168 (N1502, N880);
nand NAND2_169 (N1505, N702, N1250);
and AND4_170 (N1507, N1251, N1252, N1253, N1254);
and AND4_171 (N1508, N1255, N1256, N1257, N1258);
nand NAND2_172 (N1509, N929, N1259);
nand NAND2_173 (N1510, N926, N1260);
nand NAND2_174 (N1511, N935, N1261);
nand NAND2_175 (N1512, N932, N1262);
and AND2_176 (N1520, N655, N1263);
and AND2_177 (N1562, N874, N1337);
not NOT1_178 (N1579, N1117);
and AND2_179 (N1580, N803, N1117);
and AND2_180 (N1581, N1338, N1345);
not NOT1_181 (N1582, N1117);
and AND2_182 (N1583, N803, N1117);
not NOT1_183 (N1584, N1117);
and AND2_184 (N1585, N803, N1117);
and AND2_185 (N1586, N854, N1347);
not NOT1_186 (N1587, N1117);
and AND2_187 (N1588, N803, N1117);
and AND2_188 (N1589, N77, N1348);
not NOT1_189 (N1590, N1117);
and AND2_190 (N1591, N803, N1117);
and AND2_191 (N1592, N1343, N1349);
not NOT1_192 (N1593, N1117);
and AND2_193 (N1594, N803, N1117);
not NOT1_194 (N1595, N1117);
and AND2_195 (N1596, N803, N1117);
and AND2_196 (N1597, N870, N1351);
not NOT1_197 (N1598, N1117);
and AND2_198 (N1599, N803, N1117);
and AND2_199 (N1600, N116, N1352);
and AND2_200 (N1643, N222, N1401);
and AND2_201 (N1644, N223, N1402);
and AND2_202 (N1645, N226, N1403);
and AND2_203 (N1646, N232, N1404);
and AND2_204 (N1647, N238, N1405);
and AND2_205 (N1648, N244, N1406);
and AND2_206 (N1649, N250, N1407);
and AND2_207 (N1650, N257, N1408);
and AND3_208 (N1667, N1, N13, N1426);
and AND3_209 (N1670, N1, N13, N1427);
not NOT1_210 (N1673, N1202);
not NOT1_211 (N1674, N1202);
not NOT1_212 (N1675, N1202);
not NOT1_213 (N1676, N1202);
not NOT1_214 (N1677, N1202);
not NOT1_215 (N1678, N1202);
not NOT1_216 (N1679, N1202);
not NOT1_217 (N1680, N1202);
nand NAND2_218 (N1691, N941, N1467);
nand NAND2_219 (N1692, N938, N1468);
nand NAND2_220 (N1693, N947, N1469);
nand NAND2_221 (N1694, N944, N1470);
not NOT1_222 (N1713, N1505);
and AND2_223 (N1714, N87, N1264);
nand NAND2_224 (N1715, N1509, N1510);
nand NAND2_225 (N1718, N1511, N1512);
nand NAND2_226 (N1721, N1507, N1508);
and AND2_227 (N1722, N763, N1340);
nand NAND2_228 (N1725, N763, N1340);
not NOT1_229 (N1726, N1268);
nand NAND2_230 (N1727, N1493, N1271);
not NOT1_231 (N1728, N1493);
and AND2_232 (N1729, N683, N1268);
nand NAND2_233 (N1730, N1499, N1272);
not NOT1_234 (N1731, N1499);
nand NAND2_235 (N1735, N87, N1264);
not NOT1_236 (N1736, N1273);
not NOT1_237 (N1737, N1276);
nand NAND2_238 (N1738, N1325, N821);
nand NAND2_239 (N1747, N1325, N825);
nand NAND3_240 (N1756, N772, N1279, N798);
nand NAND4_241 (N1761, N772, N786, N798, N1302);
nand NAND2_242 (N1764, N1496, N1339);
not NOT1_243 (N1765, N1496);
nand NAND2_244 (N1766, N1502, N1344);
not NOT1_245 (N1767, N1502);
not NOT1_246 (N1768, N1328);
not NOT1_247 (N1769, N1334);
not NOT1_248 (N1770, N1331);
and AND2_249 (N1787, N845, N1579);
and AND2_250 (N1788, N150, N1580);
and AND2_251 (N1789, N851, N1582);
and AND2_252 (N1790, N159, N1583);
and AND2_253 (N1791, N77, N1584);
and AND2_254 (N1792, N50, N1585);
and AND2_255 (N1793, N858, N1587);
and AND2_256 (N1794, N845, N1588);
and AND2_257 (N1795, N864, N1590);
and AND2_258 (N1796, N851, N1591);
and AND2_259 (N1797, N107, N1593);
and AND2_260 (N1798, N77, N1594);
and AND2_261 (N1799, N116, N1595);
and AND2_262 (N1800, N858, N1596);
and AND2_263 (N1801, N283, N1598);
and AND2_264 (N1802, N864, N1599);
and AND2_265 (N1803, N200, N1363);
and AND2_266 (N1806, N889, N1363);
and AND2_267 (N1809, N890, N1366);
and AND2_268 (N1812, N891, N1366);
nand NAND2_269 (N1815, N1298, N1302);
nand NAND2_270 (N1818, N821, N1302);
nand NAND3_271 (N1821, N772, N1279, N1179);
nand NAND3_272 (N1824, N786, N794, N1298);
nand NAND2_273 (N1833, N786, N1298);
not NOT1_274 (N1842, N1369);
not NOT1_275 (N1843, N1369);
not NOT1_276 (N1844, N1369);
not NOT1_277 (N1845, N1369);
not NOT1_278 (N1846, N1369);
not NOT1_279 (N1847, N1369);
not NOT1_280 (N1848, N1369);
not NOT1_281 (N1849, N1384);
and AND2_282 (N1850, N1384, N896);
not NOT1_283 (N1851, N1384);
and AND2_284 (N1852, N1384, N896);
not NOT1_285 (N1853, N1384);
and AND2_286 (N1854, N1384, N896);
not NOT1_287 (N1855, N1384);
and AND2_288 (N1856, N1384, N896);
not NOT1_289 (N1857, N1384);
and AND2_290 (N1858, N1384, N896);
not NOT1_291 (N1859, N1384);
and AND2_292 (N1860, N1384, N896);
not NOT1_293 (N1861, N1384);
and AND2_294 (N1862, N1384, N896);
not NOT1_295 (N1863, N1384);
and AND2_296 (N1864, N1384, N896);
and AND2_297 (N1869, N1202, N1409);
nor NOR2_298 (N1870, N50, N1409);
not NOT1_299 (N1873, N1306);
and AND2_300 (N1874, N1202, N1409);
nor NOR2_301 (N1875, N58, N1409);
not NOT1_302 (N1878, N1306);
and AND2_303 (N1879, N1202, N1409);
nor NOR2_304 (N1880, N68, N1409);
not NOT1_305 (N1883, N1306);
and AND2_306 (N1884, N1202, N1409);
nor NOR2_307 (N1885, N77, N1409);
not NOT1_308 (N1888, N1306);
and AND2_309 (N1889, N1202, N1409);
nor NOR2_310 (N1890, N87, N1409);
not NOT1_311 (N1893, N1322);
and AND2_312 (N1894, N1202, N1409);
nor NOR2_313 (N1895, N97, N1409);
not NOT1_314 (N1898, N1315);
and AND2_315 (N1899, N1202, N1409);
nor NOR2_316 (N1900, N107, N1409);
not NOT1_317 (N1903, N1315);
and AND2_318 (N1904, N1202, N1409);
nor NOR2_319 (N1905, N116, N1409);
not NOT1_320 (N1908, N1315);
and AND2_321 (N1909, N1452, N213);
nand NAND2_322 (N1912, N1452, N213);
and AND3_323 (N1913, N1452, N213, N343);
nand NAND3_324 (N1917, N1452, N213, N343);
and AND3_325 (N1922, N1452, N213, N343);
nand NAND3_326 (N1926, N1452, N213, N343);
buf BUFF1_327 (N1930, N1464);
nand NAND2_328 (N1933, N1691, N1692);
nand NAND2_329 (N1936, N1693, N1694);
not NOT1_330 (N1939, N1471);
nand NAND2_331 (N1940, N1471, N1474);
not NOT1_332 (N1941, N1475);
not NOT1_333 (N1942, N1478);
not NOT1_334 (N1943, N1481);
not NOT1_335 (N1944, N1484);
not NOT1_336 (N1945, N1487);
not NOT1_337 (N1946, N1490);
not NOT1_338 (N1947, N1714);
nand NAND2_339 (N1960, N953, N1728);
nand NAND2_340 (N1961, N959, N1731);
and AND2_341 (N1966, N1520, N1276);
nand NAND2_342 (N1981, N956, N1765);
nand NAND2_343 (N1982, N962, N1767);
and AND2_344 (N1983, N1067, N1768);
or OR3_345 (N1986, N1581, N1787, N1788);
or OR3_346 (N1987, N1586, N1791, N1792);
or OR3_347 (N1988, N1589, N1793, N1794);
or OR3_348 (N1989, N1592, N1795, N1796);
or OR3_349 (N1990, N1597, N1799, N1800);
or OR3_350 (N1991, N1600, N1801, N1802);
and AND2_351 (N2022, N77, N1849);
and AND2_352 (N2023, N223, N1850);
and AND2_353 (N2024, N87, N1851);
and AND2_354 (N2025, N226, N1852);
and AND2_355 (N2026, N97, N1853);
and AND2_356 (N2027, N232, N1854);
and AND2_357 (N2028, N107, N1855);
and AND2_358 (N2029, N238, N1856);
and AND2_359 (N2030, N116, N1857);
and AND2_360 (N2031, N244, N1858);
and AND2_361 (N2032, N283, N1859);
and AND2_362 (N2033, N250, N1860);
and AND2_363 (N2034, N294, N1861);
and AND2_364 (N2035, N257, N1862);
and AND2_365 (N2036, N303, N1863);
and AND2_366 (N2037, N264, N1864);
buf BUFF1_367 (N2038, N1667);
not NOT1_368 (N2043, N1667);
buf BUFF1_369 (N2052, N1670);
not NOT1_370 (N2057, N1670);
and AND3_371 (N2068, N50, N1197, N1869);
and AND3_372 (N2073, N58, N1197, N1874);
and AND3_373 (N2078, N68, N1197, N1879);
and AND3_374 (N2083, N77, N1197, N1884);
and AND3_375 (N2088, N87, N1219, N1889);
and AND3_376 (N2093, N97, N1219, N1894);
and AND3_377 (N2098, N107, N1219, N1899);
and AND3_378 (N2103, N116, N1219, N1904);
not NOT1_379 (N2121, N1562);
not NOT1_380 (N2122, N1562);
not NOT1_381 (N2123, N1562);
not NOT1_382 (N2124, N1562);
not NOT1_383 (N2125, N1562);
not NOT1_384 (N2126, N1562);
not NOT1_385 (N2127, N1562);
not NOT1_386 (N2128, N1562);
nand NAND2_387 (N2133, N950, N1939);
nand NAND2_388 (N2134, N1478, N1941);
nand NAND2_389 (N2135, N1475, N1942);
nand NAND2_390 (N2136, N1484, N1943);
nand NAND2_391 (N2137, N1481, N1944);
nand NAND2_392 (N2138, N1490, N1945);
nand NAND2_393 (N2139, N1487, N1946);
not NOT1_394 (N2141, N1933);
not NOT1_395 (N2142, N1936);
not NOT1_396 (N2143, N1738);
and AND2_397 (N2144, N1738, N1747);
not NOT1_398 (N2145, N1747);
nand NAND2_399 (N2146, N1727, N1960);
nand NAND2_400 (N2147, N1730, N1961);
and AND4_401 (N2148, N1722, N1267, N665, N58);
not NOT1_402 (N2149, N1738);
and AND2_403 (N2150, N1738, N1747);
not NOT1_404 (N2151, N1747);
not NOT1_405 (N2152, N1738);
not NOT1_406 (N2153, N1747);
and AND2_407 (N2154, N1738, N1747);
not NOT1_408 (N2155, N1738);
not NOT1_409 (N2156, N1747);
and AND2_410 (N2157, N1738, N1747);
buf BUFF1_411 (N2158, N1761);
buf BUFF1_412 (N2175, N1761);
nand NAND2_413 (N2178, N1764, N1981);
nand NAND2_414 (N2179, N1766, N1982);
not NOT1_415 (N2180, N1756);
and AND2_416 (N2181, N1756, N1328);
not NOT1_417 (N2183, N1756);
and AND2_418 (N2184, N1331, N1756);
nand NAND2_419 (N2185, N1358, N1812);
nand NAND2_420 (N2188, N1358, N1809);
nand NAND2_421 (N2191, N1353, N1812);
nand NAND2_422 (N2194, N1353, N1809);
nand NAND2_423 (N2197, N1358, N1806);
nand NAND2_424 (N2200, N1358, N1803);
nand NAND2_425 (N2203, N1353, N1806);
nand NAND2_426 (N2206, N1353, N1803);
not NOT1_427 (N2209, N1815);
not NOT1_428 (N2210, N1818);
and AND2_429 (N2211, N1815, N1818);
buf BUFF1_430 (N2212, N1821);
buf BUFF1_431 (N2221, N1821);
not NOT1_432 (N2230, N1833);
not NOT1_433 (N2231, N1833);
not NOT1_434 (N2232, N1833);
not NOT1_435 (N2233, N1833);
not NOT1_436 (N2234, N1824);
not NOT1_437 (N2235, N1824);
not NOT1_438 (N2236, N1824);
not NOT1_439 (N2237, N1824);
or OR3_440 (N2238, N2022, N1643, N2023);
or OR3_441 (N2239, N2024, N1644, N2025);
or OR3_442 (N2240, N2026, N1645, N2027);
or OR3_443 (N2241, N2028, N1646, N2029);
or OR3_444 (N2242, N2030, N1647, N2031);
or OR3_445 (N2243, N2032, N1648, N2033);
or OR3_446 (N2244, N2034, N1649, N2035);
or OR3_447 (N2245, N2036, N1650, N2037);
and AND2_448 (N2270, N1986, N1673);
and AND2_449 (N2277, N1987, N1675);
and AND2_450 (N2282, N1988, N1676);
and AND2_451 (N2287, N1989, N1677);
and AND2_452 (N2294, N1990, N1679);
and AND2_453 (N2299, N1991, N1680);
buf BUFF1_454 (N2304, N1917);
and AND2_455 (N2307, N1930, N350);
nand NAND2_456 (N2310, N1930, N350);
buf BUFF1_457 (N2313, N1715);
buf BUFF1_458 (N2316, N1718);
buf BUFF1_459 (N2319, N1715);
buf BUFF1_460 (N2322, N1718);
nand NAND2_461 (N2325, N1940, N2133);
nand NAND2_462 (N2328, N2134, N2135);
nand NAND2_463 (N2331, N2136, N2137);
nand NAND2_464 (N2334, N2138, N2139);
nand NAND2_465 (N2341, N1936, N2141);
nand NAND2_466 (N2342, N1933, N2142);
and AND2_467 (N2347, N724, N2144);
and AND3_468 (N2348, N2146, N699, N1726);
and AND2_469 (N2349, N753, N2147);
and AND2_470 (N2350, N2148, N1273);
and AND2_471 (N2351, N736, N2150);
and AND2_472 (N2352, N1735, N2153);
and AND2_473 (N2353, N763, N2154);
and AND2_474 (N2354, N1725, N2156);
and AND2_475 (N2355, N749, N2157);
not NOT1_476 (N2374, N2178);
not NOT1_477 (N2375, N2179);
and AND2_478 (N2376, N1520, N2180);
and AND2_479 (N2379, N1721, N2181);
and AND2_480 (N2398, N665, N2211);
and AND3_481 (N2417, N2057, N226, N1873);
and AND3_482 (N2418, N2057, N274, N1306);
and AND2_483 (N2419, N2052, N2238);
and AND3_484 (N2420, N2057, N232, N1878);
and AND3_485 (N2421, N2057, N274, N1306);
and AND2_486 (N2422, N2052, N2239);
and AND3_487 (N2425, N2057, N238, N1883);
and AND3_488 (N2426, N2057, N274, N1306);
and AND2_489 (N2427, N2052, N2240);
and AND3_490 (N2430, N2057, N244, N1888);
and AND3_491 (N2431, N2057, N274, N1306);
and AND2_492 (N2432, N2052, N2241);
and AND3_493 (N2435, N2043, N250, N1893);
and AND3_494 (N2436, N2043, N274, N1322);
and AND2_495 (N2437, N2038, N2242);
and AND3_496 (N2438, N2043, N257, N1898);
and AND3_497 (N2439, N2043, N274, N1315);
and AND2_498 (N2440, N2038, N2243);
and AND3_499 (N2443, N2043, N264, N1903);
and AND3_500 (N2444, N2043, N274, N1315);
and AND2_501 (N2445, N2038, N2244);
and AND3_502 (N2448, N2043, N270, N1908);
and AND3_503 (N2449, N2043, N274, N1315);
and AND2_504 (N2450, N2038, N2245);
not NOT1_505 (N2467, N2313);
not NOT1_506 (N2468, N2316);
not NOT1_507 (N2469, N2319);
not NOT1_508 (N2470, N2322);
nand NAND2_509 (N2471, N2341, N2342);
not NOT1_510 (N2474, N2325);
not NOT1_511 (N2475, N2328);
not NOT1_512 (N2476, N2331);
not NOT1_513 (N2477, N2334);
or OR2_514 (N2478, N2348, N1729);
not NOT1_515 (N2481, N2175);
and AND2_516 (N2482, N2175, N1334);
and AND2_517 (N2483, N2349, N2183);
and AND2_518 (N2486, N2374, N1346);
and AND2_519 (N2487, N2375, N1350);
buf BUFF1_520 (N2488, N2185);
buf BUFF1_521 (N2497, N2188);
buf BUFF1_522 (N2506, N2191);
buf BUFF1_523 (N2515, N2194);
buf BUFF1_524 (N2524, N2197);
buf BUFF1_525 (N2533, N2200);
buf BUFF1_526 (N2542, N2203);
buf BUFF1_527 (N2551, N2206);
buf BUFF1_528 (N2560, N2185);
buf BUFF1_529 (N2569, N2188);
buf BUFF1_530 (N2578, N2191);
buf BUFF1_531 (N2587, N2194);
buf BUFF1_532 (N2596, N2197);
buf BUFF1_533 (N2605, N2200);
buf BUFF1_534 (N2614, N2203);
buf BUFF1_535 (N2623, N2206);
not NOT1_536 (N2632, N2212);
and AND2_537 (N2633, N2212, N1833);
not NOT1_538 (N2634, N2212);
and AND2_539 (N2635, N2212, N1833);
not NOT1_540 (N2636, N2212);
and AND2_541 (N2637, N2212, N1833);
not NOT1_542 (N2638, N2212);
and AND2_543 (N2639, N2212, N1833);
not NOT1_544 (N2640, N2221);
and AND2_545 (N2641, N2221, N1824);
not NOT1_546 (N2642, N2221);
and AND2_547 (N2643, N2221, N1824);
not NOT1_548 (N2644, N2221);
and AND2_549 (N2645, N2221, N1824);
not NOT1_550 (N2646, N2221);
and AND2_551 (N2647, N2221, N1824);
or OR3_552 (N2648, N2270, N1870, N2068);
nor NOR3_553 (N2652, N2270, N1870, N2068);
or OR3_554 (N2656, N2417, N2418, N2419);
or OR3_555 (N2659, N2420, N2421, N2422);
or OR3_556 (N2662, N2277, N1880, N2078);
nor NOR3_557 (N2666, N2277, N1880, N2078);
or OR3_558 (N2670, N2425, N2426, N2427);
or OR3_559 (N2673, N2282, N1885, N2083);
nor NOR3_560 (N2677, N2282, N1885, N2083);
or OR3_561 (N2681, N2430, N2431, N2432);
or OR3_562 (N2684, N2287, N1890, N2088);
nor NOR3_563 (N2688, N2287, N1890, N2088);
or OR3_564 (N2692, N2435, N2436, N2437);
or OR3_565 (N2697, N2438, N2439, N2440);
or OR3_566 (N2702, N2294, N1900, N2098);
nor NOR3_567 (N2706, N2294, N1900, N2098);
or OR3_568 (N2710, N2443, N2444, N2445);
or OR3_569 (N2715, N2299, N1905, N2103);
nor NOR3_570 (N2719, N2299, N1905, N2103);
or OR3_571 (N2723, N2448, N2449, N2450);
not NOT1_572 (N2728, N2304);
not NOT1_573 (N2729, N2158);
and AND2_574 (N2730, N1562, N2158);
not NOT1_575 (N2731, N2158);
and AND2_576 (N2732, N1562, N2158);
not NOT1_577 (N2733, N2158);
and AND2_578 (N2734, N1562, N2158);
not NOT1_579 (N2735, N2158);
and AND2_580 (N2736, N1562, N2158);
not NOT1_581 (N2737, N2158);
and AND2_582 (N2738, N1562, N2158);
not NOT1_583 (N2739, N2158);
and AND2_584 (N2740, N1562, N2158);
not NOT1_585 (N2741, N2158);
and AND2_586 (N2742, N1562, N2158);
not NOT1_587 (N2743, N2158);
and AND2_588 (N2744, N1562, N2158);
or OR3_589 (N2745, N2376, N1983, N2379);
nor NOR3_590 (N2746, N2376, N1983, N2379);
nand NAND2_591 (N2748, N2316, N2467);
nand NAND2_592 (N2749, N2313, N2468);
nand NAND2_593 (N2750, N2322, N2469);
nand NAND2_594 (N2751, N2319, N2470);
nand NAND2_595 (N2754, N2328, N2474);
nand NAND2_596 (N2755, N2325, N2475);
nand NAND2_597 (N2756, N2334, N2476);
nand NAND2_598 (N2757, N2331, N2477);
and AND2_599 (N2758, N1520, N2481);
and AND2_600 (N2761, N1722, N2482);
and AND2_601 (N2764, N2478, N1770);
or OR3_602 (N2768, N2486, N1789, N1790);
or OR3_603 (N2769, N2487, N1797, N1798);
and AND2_604 (N2898, N665, N2633);
and AND2_605 (N2899, N679, N2635);
and AND2_606 (N2900, N686, N2637);
and AND2_607 (N2901, N702, N2639);
not NOT1_608 (N2962, N2746);
nand NAND2_609 (N2966, N2748, N2749);
nand NAND2_610 (N2967, N2750, N2751);
buf BUFF1_611 (N2970, N2471);
nand NAND2_612 (N2973, N2754, N2755);
nand NAND2_613 (N2977, N2756, N2757);
and AND2_614 (N2980, N2471, N2143);
not NOT1_615 (N2984, N2488);
not NOT1_616 (N2985, N2497);
not NOT1_617 (N2986, N2506);
not NOT1_618 (N2987, N2515);
not NOT1_619 (N2988, N2524);
not NOT1_620 (N2989, N2533);
not NOT1_621 (N2990, N2542);
not NOT1_622 (N2991, N2551);
not NOT1_623 (N2992, N2488);
not NOT1_624 (N2993, N2497);
not NOT1_625 (N2994, N2506);
not NOT1_626 (N2995, N2515);
not NOT1_627 (N2996, N2524);
not NOT1_628 (N2997, N2533);
not NOT1_629 (N2998, N2542);
not NOT1_630 (N2999, N2551);
not NOT1_631 (N3000, N2488);
not NOT1_632 (N3001, N2497);
not NOT1_633 (N3002, N2506);
not NOT1_634 (N3003, N2515);
not NOT1_635 (N3004, N2524);
not NOT1_636 (N3005, N2533);
not NOT1_637 (N3006, N2542);
not NOT1_638 (N3007, N2551);
not NOT1_639 (N3008, N2488);
not NOT1_640 (N3009, N2497);
not NOT1_641 (N3010, N2506);
not NOT1_642 (N3011, N2515);
not NOT1_643 (N3012, N2524);
not NOT1_644 (N3013, N2533);
not NOT1_645 (N3014, N2542);
not NOT1_646 (N3015, N2551);
not NOT1_647 (N3016, N2488);
not NOT1_648 (N3017, N2497);
not NOT1_649 (N3018, N2506);
not NOT1_650 (N3019, N2515);
not NOT1_651 (N3020, N2524);
not NOT1_652 (N3021, N2533);
not NOT1_653 (N3022, N2542);
not NOT1_654 (N3023, N2551);
not NOT1_655 (N3024, N2488);
not NOT1_656 (N3025, N2497);
not NOT1_657 (N3026, N2506);
not NOT1_658 (N3027, N2515);
not NOT1_659 (N3028, N2524);
not NOT1_660 (N3029, N2533);
not NOT1_661 (N3030, N2542);
not NOT1_662 (N3031, N2551);
not NOT1_663 (N3032, N2488);
not NOT1_664 (N3033, N2497);
not NOT1_665 (N3034, N2506);
not NOT1_666 (N3035, N2515);
not NOT1_667 (N3036, N2524);
not NOT1_668 (N3037, N2533);
not NOT1_669 (N3038, N2542);
not NOT1_670 (N3039, N2551);
not NOT1_671 (N3040, N2488);
not NOT1_672 (N3041, N2497);
not NOT1_673 (N3042, N2506);
not NOT1_674 (N3043, N2515);
not NOT1_675 (N3044, N2524);
not NOT1_676 (N3045, N2533);
not NOT1_677 (N3046, N2542);
not NOT1_678 (N3047, N2551);
not NOT1_679 (N3048, N2560);
not NOT1_680 (N3049, N2569);
not NOT1_681 (N3050, N2578);
not NOT1_682 (N3051, N2587);
not NOT1_683 (N3052, N2596);
not NOT1_684 (N3053, N2605);
not NOT1_685 (N3054, N2614);
not NOT1_686 (N3055, N2623);
not NOT1_687 (N3056, N2560);
not NOT1_688 (N3057, N2569);
not NOT1_689 (N3058, N2578);
not NOT1_690 (N3059, N2587);
not NOT1_691 (N3060, N2596);
not NOT1_692 (N3061, N2605);
not NOT1_693 (N3062, N2614);
not NOT1_694 (N3063, N2623);
not NOT1_695 (N3064, N2560);
not NOT1_696 (N3065, N2569);
not NOT1_697 (N3066, N2578);
not NOT1_698 (N3067, N2587);
not NOT1_699 (N3068, N2596);
not NOT1_700 (N3069, N2605);
not NOT1_701 (N3070, N2614);
not NOT1_702 (N3071, N2623);
not NOT1_703 (N3072, N2560);
not NOT1_704 (N3073, N2569);
not NOT1_705 (N3074, N2578);
not NOT1_706 (N3075, N2587);
not NOT1_707 (N3076, N2596);
not NOT1_708 (N3077, N2605);
not NOT1_709 (N3078, N2614);
not NOT1_710 (N3079, N2623);
not NOT1_711 (N3080, N2560);
not NOT1_712 (N3081, N2569);
not NOT1_713 (N3082, N2578);
not NOT1_714 (N3083, N2587);
not NOT1_715 (N3084, N2596);
not NOT1_716 (N3085, N2605);
not NOT1_717 (N3086, N2614);
not NOT1_718 (N3087, N2623);
not NOT1_719 (N3088, N2560);
not NOT1_720 (N3089, N2569);
not NOT1_721 (N3090, N2578);
not NOT1_722 (N3091, N2587);
not NOT1_723 (N3092, N2596);
not NOT1_724 (N3093, N2605);
not NOT1_725 (N3094, N2614);
not NOT1_726 (N3095, N2623);
not NOT1_727 (N3096, N2560);
not NOT1_728 (N3097, N2569);
not NOT1_729 (N3098, N2578);
not NOT1_730 (N3099, N2587);
not NOT1_731 (N3100, N2596);
not NOT1_732 (N3101, N2605);
not NOT1_733 (N3102, N2614);
not NOT1_734 (N3103, N2623);
not NOT1_735 (N3104, N2560);
not NOT1_736 (N3105, N2569);
not NOT1_737 (N3106, N2578);
not NOT1_738 (N3107, N2587);
not NOT1_739 (N3108, N2596);
not NOT1_740 (N3109, N2605);
not NOT1_741 (N3110, N2614);
not NOT1_742 (N3111, N2623);
buf BUFF1_743 (N3112, N2656);
not NOT1_744 (N3115, N2656);
not NOT1_745 (N3118, N2652);
and AND2_746 (N3119, N2768, N1674);
buf BUFF1_747 (N3122, N2659);
not NOT1_748 (N3125, N2659);
buf BUFF1_749 (N3128, N2670);
not NOT1_750 (N3131, N2670);
not NOT1_751 (N3134, N2666);
buf BUFF1_752 (N3135, N2681);
not NOT1_753 (N3138, N2681);
not NOT1_754 (N3141, N2677);
buf BUFF1_755 (N3142, N2692);
not NOT1_756 (N3145, N2692);
not NOT1_757 (N3148, N2688);
and AND2_758 (N3149, N2769, N1678);
buf BUFF1_759 (N3152, N2697);
not NOT1_760 (N3155, N2697);
buf BUFF1_761 (N3158, N2710);
not NOT1_762 (N3161, N2710);
not NOT1_763 (N3164, N2706);
buf BUFF1_764 (N3165, N2723);
not NOT1_765 (N3168, N2723);
not NOT1_766 (N3171, N2719);
and AND2_767 (N3172, N1909, N2648);
and AND2_768 (N3175, N1913, N2662);
and AND2_769 (N3178, N1913, N2673);
and AND2_770 (N3181, N1913, N2684);
and AND2_771 (N3184, N1922, N2702);
and AND2_772 (N3187, N1922, N2715);
not NOT1_773 (N3190, N2692);
not NOT1_774 (N3191, N2697);
not NOT1_775 (N3192, N2710);
not NOT1_776 (N3193, N2723);
and AND5_777 (N3194, N2692, N2697, N2710, N2723, N1459);
nand NAND2_778 (N3195, N2745, N2962);
not NOT1_779 (N3196, N2966);
or OR3_780 (N3206, N2980, N2145, N2347);
and AND2_781 (N3207, N124, N2984);
and AND2_782 (N3208, N159, N2985);
and AND2_783 (N3209, N150, N2986);
and AND2_784 (N3210, N143, N2987);
and AND2_785 (N3211, N137, N2988);
and AND2_786 (N3212, N132, N2989);
and AND2_787 (N3213, N128, N2990);
and AND2_788 (N3214, N125, N2991);
and AND2_789 (N3215, N125, N2992);
and AND2_790 (N3216, N655, N2993);
and AND2_791 (N3217, N159, N2994);
and AND2_792 (N3218, N150, N2995);
and AND2_793 (N3219, N143, N2996);
and AND2_794 (N3220, N137, N2997);
and AND2_795 (N3221, N132, N2998);
and AND2_796 (N3222, N128, N2999);
and AND2_797 (N3223, N128, N3000);
and AND2_798 (N3224, N670, N3001);
and AND2_799 (N3225, N655, N3002);
and AND2_800 (N3226, N159, N3003);
and AND2_801 (N3227, N150, N3004);
and AND2_802 (N3228, N143, N3005);
and AND2_803 (N3229, N137, N3006);
and AND2_804 (N3230, N132, N3007);
and AND2_805 (N3231, N132, N3008);
and AND2_806 (N3232, N690, N3009);
and AND2_807 (N3233, N670, N3010);
and AND2_808 (N3234, N655, N3011);
and AND2_809 (N3235, N159, N3012);
and AND2_810 (N3236, N150, N3013);
and AND2_811 (N3237, N143, N3014);
and AND2_812 (N3238, N137, N3015);
and AND2_813 (N3239, N137, N3016);
and AND2_814 (N3240, N706, N3017);
and AND2_815 (N3241, N690, N3018);
and AND2_816 (N3242, N670, N3019);
and AND2_817 (N3243, N655, N3020);
and AND2_818 (N3244, N159, N3021);
and AND2_819 (N3245, N150, N3022);
and AND2_820 (N3246, N143, N3023);
and AND2_821 (N3247, N143, N3024);
and AND2_822 (N3248, N715, N3025);
and AND2_823 (N3249, N706, N3026);
and AND2_824 (N3250, N690, N3027);
and AND2_825 (N3251, N670, N3028);
and AND2_826 (N3252, N655, N3029);
and AND2_827 (N3253, N159, N3030);
and AND2_828 (N3254, N150, N3031);
and AND2_829 (N3255, N150, N3032);
and AND2_830 (N3256, N727, N3033);
and AND2_831 (N3257, N715, N3034);
and AND2_832 (N3258, N706, N3035);
and AND2_833 (N3259, N690, N3036);
and AND2_834 (N3260, N670, N3037);
and AND2_835 (N3261, N655, N3038);
and AND2_836 (N3262, N159, N3039);
and AND2_837 (N3263, N159, N3040);
and AND2_838 (N3264, N740, N3041);
and AND2_839 (N3265, N727, N3042);
and AND2_840 (N3266, N715, N3043);
and AND2_841 (N3267, N706, N3044);
and AND2_842 (N3268, N690, N3045);
and AND2_843 (N3269, N670, N3046);
and AND2_844 (N3270, N655, N3047);
and AND2_845 (N3271, N283, N3048);
and AND2_846 (N3272, N670, N3049);
and AND2_847 (N3273, N690, N3050);
and AND2_848 (N3274, N706, N3051);
and AND2_849 (N3275, N715, N3052);
and AND2_850 (N3276, N727, N3053);
and AND2_851 (N3277, N740, N3054);
and AND2_852 (N3278, N753, N3055);
and AND2_853 (N3279, N294, N3056);
and AND2_854 (N3280, N690, N3057);
and AND2_855 (N3281, N706, N3058);
and AND2_856 (N3282, N715, N3059);
and AND2_857 (N3283, N727, N3060);
and AND2_858 (N3284, N740, N3061);
and AND2_859 (N3285, N753, N3062);
and AND2_860 (N3286, N283, N3063);
and AND2_861 (N3287, N303, N3064);
and AND2_862 (N3288, N706, N3065);
and AND2_863 (N3289, N715, N3066);
and AND2_864 (N3290, N727, N3067);
and AND2_865 (N3291, N740, N3068);
and AND2_866 (N3292, N753, N3069);
and AND2_867 (N3293, N283, N3070);
and AND2_868 (N3294, N294, N3071);
and AND2_869 (N3295, N311, N3072);
and AND2_870 (N3296, N715, N3073);
and AND2_871 (N3297, N727, N3074);
and AND2_872 (N3298, N740, N3075);
and AND2_873 (N3299, N753, N3076);
and AND2_874 (N3300, N283, N3077);
and AND2_875 (N3301, N294, N3078);
and AND2_876 (N3302, N303, N3079);
and AND2_877 (N3303, N317, N3080);
and AND2_878 (N3304, N727, N3081);
and AND2_879 (N3305, N740, N3082);
and AND2_880 (N3306, N753, N3083);
and AND2_881 (N3307, N283, N3084);
and AND2_882 (N3308, N294, N3085);
and AND2_883 (N3309, N303, N3086);
and AND2_884 (N3310, N311, N3087);
and AND2_885 (N3311, N322, N3088);
and AND2_886 (N3312, N740, N3089);
and AND2_887 (N3313, N753, N3090);
and AND2_888 (N3314, N283, N3091);
and AND2_889 (N3315, N294, N3092);
and AND2_890 (N3316, N303, N3093);
and AND2_891 (N3317, N311, N3094);
and AND2_892 (N3318, N317, N3095);
and AND2_893 (N3319, N326, N3096);
and AND2_894 (N3320, N753, N3097);
and AND2_895 (N3321, N283, N3098);
and AND2_896 (N3322, N294, N3099);
and AND2_897 (N3323, N303, N3100);
and AND2_898 (N3324, N311, N3101);
and AND2_899 (N3325, N317, N3102);
and AND2_900 (N3326, N322, N3103);
and AND2_901 (N3327, N329, N3104);
and AND2_902 (N3328, N283, N3105);
and AND2_903 (N3329, N294, N3106);
and AND2_904 (N3330, N303, N3107);
and AND2_905 (N3331, N311, N3108);
and AND2_906 (N3332, N317, N3109);
and AND2_907 (N3333, N322, N3110);
and AND2_908 (N3334, N326, N3111);
and AND5_909 (N3383, N3190, N3191, N3192, N3193, N917);
buf BUFF1_910 (N3384, N2977);
and AND2_911 (N3387, N3196, N1736);
and AND2_912 (N3388, N2977, N2149);
and AND2_913 (N3389, N2973, N1737);
nor NOR8_914 (N3390, N3207, N3208, N3209, N3210, N3211, N3212, N3213, N3214);
nor NOR8_915 (N3391, N3215, N3216, N3217, N3218, N3219, N3220, N3221, N3222);
nor NOR8_916 (N3392, N3223, N3224, N3225, N3226, N3227, N3228, N3229, N3230);
nor NOR8_917 (N3393, N3231, N3232, N3233, N3234, N3235, N3236, N3237, N3238);
nor NOR8_918 (N3394, N3239, N3240, N3241, N3242, N3243, N3244, N3245, N3246);
nor NOR8_919 (N3395, N3247, N3248, N3249, N3250, N3251, N3252, N3253, N3254);
nor NOR8_920 (N3396, N3255, N3256, N3257, N3258, N3259, N3260, N3261, N3262);
nor NOR8_921 (N3397, N3263, N3264, N3265, N3266, N3267, N3268, N3269, N3270);
nor NOR8_922 (N3398, N3271, N3272, N3273, N3274, N3275, N3276, N3277, N3278);
nor NOR8_923 (N3399, N3279, N3280, N3281, N3282, N3283, N3284, N3285, N3286);
nor NOR8_924 (N3400, N3287, N3288, N3289, N3290, N3291, N3292, N3293, N3294);
nor NOR8_925 (N3401, N3295, N3296, N3297, N3298, N3299, N3300, N3301, N3302);
nor NOR8_926 (N3402, N3303, N3304, N3305, N3306, N3307, N3308, N3309, N3310);
nor NOR8_927 (N3403, N3311, N3312, N3313, N3314, N3315, N3316, N3317, N3318);
nor NOR8_928 (N3404, N3319, N3320, N3321, N3322, N3323, N3324, N3325, N3326);
nor NOR8_929 (N3405, N3327, N3328, N3329, N3330, N3331, N3332, N3333, N3334);
and AND2_930 (N3406, N3206, N2641);
and AND3_931 (N3407, N169, N2648, N3112);
and AND3_932 (N3410, N179, N2648, N3115);
and AND3_933 (N3413, N190, N2652, N3115);
and AND3_934 (N3414, N200, N2652, N3112);
or OR3_935 (N3415, N3119, N1875, N2073);
nor NOR3_936 (N3419, N3119, N1875, N2073);
and AND3_937 (N3423, N169, N2662, N3128);
and AND3_938 (N3426, N179, N2662, N3131);
and AND3_939 (N3429, N190, N2666, N3131);
and AND3_940 (N3430, N200, N2666, N3128);
and AND3_941 (N3431, N169, N2673, N3135);
and AND3_942 (N3434, N179, N2673, N3138);
and AND3_943 (N3437, N190, N2677, N3138);
and AND3_944 (N3438, N200, N2677, N3135);
and AND3_945 (N3439, N169, N2684, N3142);
and AND3_946 (N3442, N179, N2684, N3145);
and AND3_947 (N3445, N190, N2688, N3145);
and AND3_948 (N3446, N200, N2688, N3142);
or OR3_949 (N3447, N3149, N1895, N2093);
nor NOR3_950 (N3451, N3149, N1895, N2093);
and AND3_951 (N3455, N169, N2702, N3158);
and AND3_952 (N3458, N179, N2702, N3161);
and AND3_953 (N3461, N190, N2706, N3161);
and AND3_954 (N3462, N200, N2706, N3158);
and AND3_955 (N3463, N169, N2715, N3165);
and AND3_956 (N3466, N179, N2715, N3168);
and AND3_957 (N3469, N190, N2719, N3168);
and AND3_958 (N3470, N200, N2719, N3165);
or OR2_959 (N3471, N3194, N3383);
buf BUFF1_960 (N3472, N2967);
buf BUFF1_961 (N3475, N2970);
buf BUFF1_962 (N3478, N2967);
buf BUFF1_963 (N3481, N2970);
buf BUFF1_964 (N3484, N2973);
buf BUFF1_965 (N3487, N2973);
buf BUFF1_966 (N3490, N3172);
buf BUFF1_967 (N3493, N3172);
buf BUFF1_968 (N3496, N3175);
buf BUFF1_969 (N3499, N3175);
buf BUFF1_970 (N3502, N3178);
buf BUFF1_971 (N3505, N3178);
buf BUFF1_972 (N3508, N3181);
buf BUFF1_973 (N3511, N3181);
buf BUFF1_974 (N3514, N3184);
buf BUFF1_975 (N3517, N3184);
buf BUFF1_976 (N3520, N3187);
buf BUFF1_977 (N3523, N3187);
nor NOR2_978 (N3534, N3387, N2350);
or OR3_979 (N3535, N3388, N2151, N2351);
nor NOR2_980 (N3536, N3389, N1966);
and AND2_981 (N3537, N3390, N2209);
and AND2_982 (N3538, N3398, N2210);
and AND2_983 (N3539, N3391, N1842);
and AND2_984 (N3540, N3399, N1369);
and AND2_985 (N3541, N3392, N1843);
and AND2_986 (N3542, N3400, N1369);
and AND2_987 (N3543, N3393, N1844);
and AND2_988 (N3544, N3401, N1369);
and AND2_989 (N3545, N3394, N1845);
and AND2_990 (N3546, N3402, N1369);
and AND2_991 (N3547, N3395, N1846);
and AND2_992 (N3548, N3403, N1369);
and AND2_993 (N3549, N3396, N1847);
and AND2_994 (N3550, N3404, N1369);
and AND2_995 (N3551, N3397, N1848);
and AND2_996 (N3552, N3405, N1369);
or OR3_997 (N3557, N3413, N3414, N3118);
or OR3_998 (N3568, N3429, N3430, N3134);
or OR3_999 (N3573, N3437, N3438, N3141);
or OR3_1000 (N3578, N3445, N3446, N3148);
or OR3_1001 (N3589, N3461, N3462, N3164);
or OR3_1002 (N3594, N3469, N3470, N3171);
and AND2_1003 (N3605, N3471, N2728);
not NOT1_1004 (N3626, N3478);
not NOT1_1005 (N3627, N3481);
not NOT1_1006 (N3628, N3487);
not NOT1_1007 (N3629, N3484);
not NOT1_1008 (N3630, N3472);
not NOT1_1009 (N3631, N3475);
and AND2_1010 (N3632, N3536, N2152);
and AND2_1011 (N3633, N3534, N2155);
or OR3_1012 (N3634, N3537, N3538, N2398);
or OR2_1013 (N3635, N3539, N3540);
or OR2_1014 (N3636, N3541, N3542);
or OR2_1015 (N3637, N3543, N3544);
or OR2_1016 (N3638, N3545, N3546);
or OR2_1017 (N3639, N3547, N3548);
or OR2_1018 (N3640, N3549, N3550);
or OR2_1019 (N3641, N3551, N3552);
and AND2_1020 (N3642, N3535, N2643);
or OR2_1021 (N3643, N3407, N3410);
nor NOR2_1022 (N3644, N3407, N3410);
and AND3_1023 (N3645, N169, N3415, N3122);
and AND3_1024 (N3648, N179, N3415, N3125);
and AND3_1025 (N3651, N190, N3419, N3125);
and AND3_1026 (N3652, N200, N3419, N3122);
not NOT1_1027 (N3653, N3419);
or OR2_1028 (N3654, N3423, N3426);
nor NOR2_1029 (N3657, N3423, N3426);
or OR2_1030 (N3658, N3431, N3434);
nor NOR2_1031 (N3661, N3431, N3434);
or OR2_1032 (N3662, N3439, N3442);
nor NOR2_1033 (N3663, N3439, N3442);
and AND3_1034 (N3664, N169, N3447, N3152);
and AND3_1035 (N3667, N179, N3447, N3155);
and AND3_1036 (N3670, N190, N3451, N3155);
and AND3_1037 (N3671, N200, N3451, N3152);
not NOT1_1038 (N3672, N3451);
or OR2_1039 (N3673, N3455, N3458);
nor NOR2_1040 (N3676, N3455, N3458);
or OR2_1041 (N3677, N3463, N3466);
nor NOR2_1042 (N3680, N3463, N3466);
not NOT1_1043 (N3681, N3493);
and AND2_1044 (N3682, N1909, N3415);
not NOT1_1045 (N3685, N3496);
not NOT1_1046 (N3686, N3499);
not NOT1_1047 (N3687, N3502);
not NOT1_1048 (N3688, N3505);
not NOT1_1049 (N3689, N3511);
and AND2_1050 (N3690, N1922, N3447);
not NOT1_1051 (N3693, N3517);
not NOT1_1052 (N3694, N3520);
not NOT1_1053 (N3695, N3523);
not NOT1_1054 (N3696, N3514);
buf BUFF1_1055 (N3697, N3384);
buf BUFF1_1056 (N3700, N3384);
not NOT1_1057 (N3703, N3490);
not NOT1_1058 (N3704, N3508);
nand NAND2_1059 (N3705, N3475, N3630);
nand NAND2_1060 (N3706, N3472, N3631);
nand NAND2_1061 (N3707, N3481, N3626);
nand NAND2_1062 (N3708, N3478, N3627);
or OR3_1063 (N3711, N3632, N2352, N2353);
or OR3_1064 (N3712, N3633, N2354, N2355);
and AND2_1065 (N3713, N3634, N2632);
and AND2_1066 (N3714, N3635, N2634);
and AND2_1067 (N3715, N3636, N2636);
and AND2_1068 (N3716, N3637, N2638);
and AND2_1069 (N3717, N3638, N2640);
and AND2_1070 (N3718, N3639, N2642);
and AND2_1071 (N3719, N3640, N2644);
and AND2_1072 (N3720, N3641, N2646);
and AND2_1073 (N3721, N3644, N3557);
or OR3_1074 (N3731, N3651, N3652, N3653);
and AND2_1075 (N3734, N3657, N3568);
and AND2_1076 (N3740, N3661, N3573);
and AND2_1077 (N3743, N3663, N3578);
or OR3_1078 (N3753, N3670, N3671, N3672);
and AND2_1079 (N3756, N3676, N3589);
and AND2_1080 (N3762, N3680, N3594);
not NOT1_1081 (N3765, N3643);
not NOT1_1082 (N3766, N3662);
nand NAND2_1083 (N3773, N3705, N3706);
nand NAND2_1084 (N3774, N3707, N3708);
nand NAND2_1085 (N3775, N3700, N3628);
not NOT1_1086 (N3776, N3700);
nand NAND2_1087 (N3777, N3697, N3629);
not NOT1_1088 (N3778, N3697);
and AND2_1089 (N3779, N3712, N2645);
and AND2_1090 (N3780, N3711, N2647);
or OR2_1091 (N3786, N3645, N3648);
nor NOR2_1092 (N3789, N3645, N3648);
or OR2_1093 (N3800, N3664, N3667);
nor NOR2_1094 (N3803, N3664, N3667);
and AND2_1095 (N3809, N3654, N1917);
and AND2_1096 (N3812, N3658, N1917);
and AND2_1097 (N3815, N3673, N1926);
and AND2_1098 (N3818, N3677, N1926);
buf BUFF1_1099 (N3821, N3682);
buf BUFF1_1100 (N3824, N3682);
buf BUFF1_1101 (N3827, N3690);
buf BUFF1_1102 (N3830, N3690);
nand NAND2_1103 (N3833, N3773, N3774);
nand NAND2_1104 (N3834, N3487, N3776);
nand NAND2_1105 (N3835, N3484, N3778);
and AND2_1106 (N3838, N3789, N3731);
and AND2_1107 (N3845, N3803, N3753);
buf BUFF1_1108 (N3850, N3721);
buf BUFF1_1109 (N3855, N3734);
buf BUFF1_1110 (N3858, N3740);
buf BUFF1_1111 (N3861, N3743);
buf BUFF1_1112 (N3865, N3756);
buf BUFF1_1113 (N3868, N3762);
nand NAND2_1114 (N3884, N3775, N3834);
nand NAND2_1115 (N3885, N3777, N3835);
nand NAND2_1116 (N3894, N3721, N3786);
nand NAND2_1117 (N3895, N3743, N3800);
not NOT1_1118 (N3898, N3821);
not NOT1_1119 (N3899, N3824);
not NOT1_1120 (N3906, N3830);
not NOT1_1121 (N3911, N3827);
and AND2_1122 (N3912, N3786, N1912);
buf BUFF1_1123 (N3913, N3812);
and AND2_1124 (N3916, N3800, N1917);
buf BUFF1_1125 (N3917, N3818);
not NOT1_1126 (N3920, N3809);
buf BUFF1_1127 (N3921, N3818);
not NOT1_1128 (N3924, N3884);
not NOT1_1129 (N3925, N3885);
and AND4_1130 (N3926, N3721, N3838, N3734, N3740);
nand NAND3_1131 (N3930, N3721, N3838, N3654);
nand NAND4_1132 (N3931, N3658, N3838, N3734, N3721);
and AND4_1133 (N3932, N3743, N3845, N3756, N3762);
nand NAND3_1134 (N3935, N3743, N3845, N3673);
nand NAND4_1135 (N3936, N3677, N3845, N3756, N3743);
buf BUFF1_1136 (N3937, N3838);
buf BUFF1_1137 (N3940, N3845);
not NOT1_1138 (N3947, N3912);
not NOT1_1139 (N3948, N3916);
buf BUFF1_1140 (N3950, N3850);
buf BUFF1_1141 (N3953, N3850);
buf BUFF1_1142 (N3956, N3855);
buf BUFF1_1143 (N3959, N3855);
buf BUFF1_1144 (N3962, N3858);
buf BUFF1_1145 (N3965, N3858);
buf BUFF1_1146 (N3968, N3861);
buf BUFF1_1147 (N3971, N3861);
buf BUFF1_1148 (N3974, N3865);
buf BUFF1_1149 (N3977, N3865);
buf BUFF1_1150 (N3980, N3868);
buf BUFF1_1151 (N3983, N3868);
nand NAND2_1152 (N3987, N3924, N3925);
nand NAND4_1153 (N3992, N3765, N3894, N3930, N3931);
nand NAND4_1154 (N3996, N3766, N3895, N3935, N3936);
not NOT1_1155 (N4013, N3921);
and AND2_1156 (N4028, N3932, N3926);
nand NAND2_1157 (N4029, N3953, N3681);
nand NAND2_1158 (N4030, N3959, N3686);
nand NAND2_1159 (N4031, N3965, N3688);
nand NAND2_1160 (N4032, N3971, N3689);
nand NAND2_1161 (N4033, N3977, N3693);
nand NAND2_1162 (N4034, N3983, N3695);
buf BUFF1_1163 (N4035, N3926);
not NOT1_1164 (N4042, N3953);
not NOT1_1165 (N4043, N3956);
nand NAND2_1166 (N4044, N3956, N3685);
not NOT1_1167 (N4045, N3959);
not NOT1_1168 (N4046, N3962);
nand NAND2_1169 (N4047, N3962, N3687);
not NOT1_1170 (N4048, N3965);
not NOT1_1171 (N4049, N3971);
not NOT1_1172 (N4050, N3977);
not NOT1_1173 (N4051, N3980);
nand NAND2_1174 (N4052, N3980, N3694);
not NOT1_1175 (N4053, N3983);
not NOT1_1176 (N4054, N3974);
nand NAND2_1177 (N4055, N3974, N3696);
and AND2_1178 (N4056, N3932, N2304);
not NOT1_1179 (N4057, N3950);
nand NAND2_1180 (N4058, N3950, N3703);
buf BUFF1_1181 (N4059, N3937);
buf BUFF1_1182 (N4062, N3937);
not NOT1_1183 (N4065, N3968);
nand NAND2_1184 (N4066, N3968, N3704);
buf BUFF1_1185 (N4067, N3940);
buf BUFF1_1186 (N4070, N3940);
nand NAND2_1187 (N4073, N3926, N3996);
not NOT1_1188 (N4074, N3992);
nand NAND2_1189 (N4075, N3493, N4042);
nand NAND2_1190 (N4076, N3499, N4045);
nand NAND2_1191 (N4077, N3505, N4048);
nand NAND2_1192 (N4078, N3511, N4049);
nand NAND2_1193 (N4079, N3517, N4050);
nand NAND2_1194 (N4080, N3523, N4053);
nand NAND2_1195 (N4085, N3496, N4043);
nand NAND2_1196 (N4086, N3502, N4046);
nand NAND2_1197 (N4088, N3520, N4051);
nand NAND2_1198 (N4090, N3514, N4054);
and AND2_1199 (N4091, N3996, N1926);
or OR2_1200 (N4094, N3605, N4056);
nand NAND2_1201 (N4098, N3490, N4057);
nand NAND2_1202 (N4101, N3508, N4065);
and AND2_1203 (N4104, N4073, N4074);
nand NAND2_1204 (N4105, N4075, N4029);
nand NAND2_1205 (N4106, N4062, N3899);
nand NAND2_1206 (N4107, N4076, N4030);
nand NAND2_1207 (N4108, N4077, N4031);
nand NAND2_1208 (N4109, N4078, N4032);
nand NAND2_1209 (N4110, N4070, N3906);
nand NAND2_1210 (N4111, N4079, N4033);
nand NAND2_1211 (N4112, N4080, N4034);
not NOT1_1212 (N4113, N4059);
nand NAND2_1213 (N4114, N4059, N3898);
not NOT1_1214 (N4115, N4062);
nand NAND2_1215 (N4116, N4085, N4044);
nand NAND2_1216 (N4119, N4086, N4047);
not NOT1_1217 (N4122, N4070);
nand NAND2_1218 (N4123, N4088, N4052);
not NOT1_1219 (N4126, N4067);
nand NAND2_1220 (N4127, N4067, N3911);
nand NAND2_1221 (N4128, N4090, N4055);
nand NAND2_1222 (N4139, N4098, N4058);
nand NAND2_1223 (N4142, N4101, N4066);
not NOT1_1224 (N4145, N4104);
not NOT1_1225 (N4146, N4105);
nand NAND2_1226 (N4147, N3824, N4115);
not NOT1_1227 (N4148, N4107);
not NOT1_1228 (N4149, N4108);
not NOT1_1229 (N4150, N4109);
nand NAND2_1230 (N4151, N3830, N4122);
not NOT1_1231 (N4152, N4111);
not NOT1_1232 (N4153, N4112);
nand NAND2_1233 (N4154, N3821, N4113);
nand NAND2_1234 (N4161, N3827, N4126);
buf BUFF1_1235 (N4167, N4091);
buf BUFF1_1236 (N4174, N4094);
buf BUFF1_1237 (N4182, N4091);
and AND2_1238 (N4186, N330, N4094);
and AND2_1239 (N4189, N4146, N2230);
nand NAND2_1240 (N4190, N4147, N4106);
and AND2_1241 (N4191, N4148, N2232);
and AND2_1242 (N4192, N4149, N2233);
and AND2_1243 (N4193, N4150, N2234);
nand NAND2_1244 (N4194, N4151, N4110);
and AND2_1245 (N4195, N4152, N2236);
and AND2_1246 (N4196, N4153, N2237);
nand NAND2_1247 (N4197, N4154, N4114);
buf BUFF1_1248 (N4200, N4116);
buf BUFF1_1249 (N4203, N4116);
buf BUFF1_1250 (N4209, N4119);
buf BUFF1_1251 (N4213, N4119);
nand NAND2_1252 (N4218, N4161, N4127);
buf BUFF1_1253 (N4223, N4123);
and AND2_1254 (N4238, N4128, N3917);
not NOT1_1255 (N4239, N4139);
not NOT1_1256 (N4241, N4142);
and AND2_1257 (N4242, N330, N4123);
buf BUFF1_1258 (N4247, N4128);
nor NOR3_1259 (N4251, N3713, N4189, N2898);
not NOT1_1260 (N4252, N4190);
nor NOR3_1261 (N4253, N3715, N4191, N2900);
nor NOR3_1262 (N4254, N3716, N4192, N2901);
nor NOR3_1263 (N4255, N3717, N4193, N3406);
not NOT1_1264 (N4256, N4194);
nor NOR3_1265 (N4257, N3719, N4195, N3779);
nor NOR3_1266 (N4258, N3720, N4196, N3780);
and AND2_1267 (N4283, N4167, N4035);
and AND2_1268 (N4284, N4174, N4035);
or OR2_1269 (N4287, N3815, N4238);
not NOT1_1270 (N4291, N4186);
not NOT1_1271 (N4295, N4167);
buf BUFF1_1272 (N4296, N4167);
not NOT1_1273 (N4299, N4182);
and AND2_1274 (N4303, N4252, N2231);
and AND2_1275 (N4304, N4256, N2235);
buf BUFF1_1276 (N4305, N4197);
or OR2_1277 (N4310, N3992, N4283);
and AND3_1278 (N4316, N4174, N4213, N4203);
and AND2_1279 (N4317, N4174, N4209);
and AND3_1280 (N4318, N4223, N4128, N4218);
and AND2_1281 (N4319, N4223, N4128);
and AND2_1282 (N4322, N4167, N4209);
nand NAND2_1283 (N4325, N4203, N3913);
nand NAND3_1284 (N4326, N4203, N4213, N4167);
nand NAND2_1285 (N4327, N4218, N3815);
nand NAND3_1286 (N4328, N4218, N4128, N3917);
nand NAND2_1287 (N4329, N4247, N4013);
not NOT1_1288 (N4330, N4247);
and AND3_1289 (N4331, N330, N4094, N4295);
and AND2_1290 (N4335, N4251, N2730);
and AND2_1291 (N4338, N4253, N2734);
and AND2_1292 (N4341, N4254, N2736);
and AND2_1293 (N4344, N4255, N2738);
and AND2_1294 (N4347, N4257, N2742);
and AND2_1295 (N4350, N4258, N2744);
buf BUFF1_1296 (N4353, N4197);
buf BUFF1_1297 (N4356, N4203);
buf BUFF1_1298 (N4359, N4209);
buf BUFF1_1299 (N4362, N4218);
buf BUFF1_1300 (N4365, N4242);
buf BUFF1_1301 (N4368, N4242);
and AND2_1302 (N4371, N4223, N4223);
nor NOR3_1303 (N4376, N3714, N4303, N2899);
nor NOR3_1304 (N4377, N3718, N4304, N3642);
and AND2_1305 (N4387, N330, N4317);
and AND2_1306 (N4390, N330, N4318);
nand NAND2_1307 (N4393, N3921, N4330);
buf BUFF1_1308 (N4398, N4287);
buf BUFF1_1309 (N4413, N4284);
nand NAND3_1310 (N4416, N3920, N4325, N4326);
or OR2_1311 (N4421, N3812, N4322);
nand NAND3_1312 (N4427, N3948, N4327, N4328);
buf BUFF1_1313 (N4430, N4287);
and AND2_1314 (N4435, N330, N4316);
or OR2_1315 (N4442, N4331, N4296);
and AND4_1316 (N4443, N4174, N4305, N4203, N4213);
nand NAND2_1317 (N4446, N4305, N3809);
nand NAND3_1318 (N4447, N4305, N4200, N3913);
nand NAND4_1319 (N4448, N4305, N4200, N4213, N4167);
not NOT1_1320 (N4452, N4356);
nand NAND2_1321 (N4458, N4329, N4393);
not NOT1_1322 (N4461, N4365);
not NOT1_1323 (N4462, N4368);
nand NAND2_1324 (N4463, N4371, N1460);
not NOT1_1325 (N4464, N4371);
buf BUFF1_1326 (N4465, N4310);
nor NOR2_1327 (N4468, N4331, N4296);
and AND2_1328 (N4472, N4376, N2732);
and AND2_1329 (N4475, N4377, N2740);
buf BUFF1_1330 (N4479, N4310);
not NOT1_1331 (N4484, N4353);
not NOT1_1332 (N4486, N4359);
nand NAND2_1333 (N4487, N4359, N4299);
not NOT1_1334 (N4491, N4362);
and AND2_1335 (N4493, N330, N4319);
not NOT1_1336 (N4496, N4398);
and AND2_1337 (N4497, N4287, N4398);
and AND2_1338 (N4498, N4442, N1769);
nand NAND4_1339 (N4503, N3947, N4446, N4447, N4448);
not NOT1_1340 (N4506, N4413);
not NOT1_1341 (N4507, N4435);
not NOT1_1342 (N4508, N4421);
nand NAND2_1343 (N4509, N4421, N4452);
not NOT1_1344 (N4510, N4427);
nand NAND2_1345 (N4511, N4427, N4241);
nand NAND2_1346 (N4515, N965, N4464);
not NOT1_1347 (N4526, N4416);
nand NAND2_1348 (N4527, N4416, N4484);
nand NAND2_1349 (N4528, N4182, N4486);
not NOT1_1350 (N4529, N4430);
nand NAND2_1351 (N4530, N4430, N4491);
buf BUFF1_1352 (N4531, N4387);
buf BUFF1_1353 (N4534, N4387);
buf BUFF1_1354 (N4537, N4390);
buf BUFF1_1355 (N4540, N4390);
and AND3_1356 (N4545, N330, N4319, N4496);
and AND2_1357 (N4549, N330, N4443);
nand NAND2_1358 (N4552, N4356, N4508);
nand NAND2_1359 (N4555, N4142, N4510);
not NOT1_1360 (N4558, N4493);
nand NAND2_1361 (N4559, N4463, N4515);
not NOT1_1362 (N4562, N4465);
and AND2_1363 (N4563, N4310, N4465);
buf BUFF1_1364 (N4564, N4468);
not NOT1_1365 (N4568, N4479);
buf BUFF1_1366 (N4569, N4443);
nand NAND2_1367 (N4572, N4353, N4526);
nand NAND2_1368 (N4573, N4362, N4529);
nand NAND2_1369 (N4576, N4487, N4528);
buf BUFF1_1370 (N4581, N4458);
buf BUFF1_1371 (N4584, N4458);
or OR3_1372 (N4587, N2758, N4498, N2761);
nor NOR3_1373 (N4588, N2758, N4498, N2761);
or OR2_1374 (N4589, N4545, N4497);
nand NAND2_1375 (N4593, N4552, N4509);
not NOT1_1376 (N4596, N4531);
not NOT1_1377 (N4597, N4534);
nand NAND2_1378 (N4599, N4555, N4511);
not NOT1_1379 (N4602, N4537);
not NOT1_1380 (N4603, N4540);
and AND3_1381 (N4608, N330, N4284, N4562);
buf BUFF1_1382 (N4613, N4503);
buf BUFF1_1383 (N4616, N4503);
nand NAND2_1384 (N4619, N4572, N4527);
nand NAND2_1385 (N4623, N4573, N4530);
not NOT1_1386 (N4628, N4588);
nand NAND2_1387 (N4629, N4569, N4506);
not NOT1_1388 (N4630, N4569);
not NOT1_1389 (N4635, N4576);
nand NAND2_1390 (N4636, N4576, N4291);
not NOT1_1391 (N4640, N4581);
nand NAND2_1392 (N4641, N4581, N4461);
not NOT1_1393 (N4642, N4584);
nand NAND2_1394 (N4643, N4584, N4462);
nor NOR2_1395 (N4644, N4608, N4563);
and AND2_1396 (N4647, N4559, N2128);
and AND2_1397 (N4650, N4559, N2743);
buf BUFF1_1398 (N4656, N4549);
buf BUFF1_1399 (N4659, N4549);
buf BUFF1_1400 (N4664, N4564);
and AND2_1401 (N4667, N4587, N4628);
nand NAND2_1402 (N4668, N4413, N4630);
not NOT1_1403 (N4669, N4616);
nand NAND2_1404 (N4670, N4616, N4239);
not NOT1_1405 (N4673, N4619);
nand NAND2_1406 (N4674, N4619, N4507);
nand NAND2_1407 (N4675, N4186, N4635);
not NOT1_1408 (N4676, N4623);
nand NAND2_1409 (N4677, N4623, N4558);
nand NAND2_1410 (N4678, N4365, N4640);
nand NAND2_1411 (N4679, N4368, N4642);
not NOT1_1412 (N4687, N4613);
nand NAND2_1413 (N4688, N4613, N4568);
buf BUFF1_1414 (N4691, N4593);
buf BUFF1_1415 (N4694, N4593);
buf BUFF1_1416 (N4697, N4599);
buf BUFF1_1417 (N4700, N4599);
nand NAND2_1418 (N4704, N4629, N4668);
nand NAND2_1419 (N4705, N4139, N4669);
not NOT1_1420 (N4706, N4656);
not NOT1_1421 (N4707, N4659);
nand NAND2_1422 (N4708, N4435, N4673);
nand NAND2_1423 (N4711, N4675, N4636);
nand NAND2_1424 (N4716, N4493, N4676);
nand NAND2_1425 (N4717, N4678, N4641);
nand NAND2_1426 (N4721, N4679, N4643);
buf BUFF1_1427 (N4722, N4644);
not NOT1_1428 (N4726, N4664);
or OR3_1429 (N4727, N4647, N4650, N4350);
nor NOR3_1430 (N4730, N4647, N4650, N4350);
nand NAND2_1431 (N4733, N4479, N4687);
nand NAND2_1432 (N4740, N4705, N4670);
nand NAND2_1433 (N4743, N4708, N4674);
not NOT1_1434 (N4747, N4691);
nand NAND2_1435 (N4748, N4691, N4596);
not NOT1_1436 (N4749, N4694);
nand NAND2_1437 (N4750, N4694, N4597);
not NOT1_1438 (N4753, N4697);
nand NAND2_1439 (N4754, N4697, N4602);
not NOT1_1440 (N4755, N4700);
nand NAND2_1441 (N4756, N4700, N4603);
nand NAND2_1442 (N4757, N4716, N4677);
nand NAND2_1443 (N4769, N4733, N4688);
and AND2_1444 (N4772, N330, N4704);
not NOT1_1445 (N4775, N4721);
not NOT1_1446 (N4778, N4730);
nand NAND2_1447 (N4786, N4531, N4747);
nand NAND2_1448 (N4787, N4534, N4749);
nand NAND2_1449 (N4788, N4537, N4753);
nand NAND2_1450 (N4789, N4540, N4755);
and AND2_1451 (N4794, N4711, N2124);
and AND2_1452 (N4797, N4711, N2735);
and AND2_1453 (N4800, N4717, N2127);
buf BUFF1_1454 (N4805, N4722);
and AND2_1455 (N4808, N4717, N4468);
buf BUFF1_1456 (N4812, N4727);
and AND2_1457 (N4815, N4727, N4778);
not NOT1_1458 (N4816, N4769);
not NOT1_1459 (N4817, N4772);
nand NAND2_1460 (N4818, N4786, N4748);
nand NAND2_1461 (N4822, N4787, N4750);
nand NAND2_1462 (N4823, N4788, N4754);
nand NAND2_1463 (N4826, N4789, N4756);
nand NAND2_1464 (N4829, N4775, N4726);
not NOT1_1465 (N4830, N4775);
and AND2_1466 (N4831, N4743, N2122);
and AND2_1467 (N4838, N4757, N2126);
buf BUFF1_1468 (N4844, N4740);
buf BUFF1_1469 (N4847, N4740);
buf BUFF1_1470 (N4850, N4743);
buf BUFF1_1471 (N4854, N4757);
nand NAND2_1472 (N4859, N4772, N4816);
nand NAND2_1473 (N4860, N4769, N4817);
not NOT1_1474 (N4868, N4826);
not NOT1_1475 (N4870, N4805);
not NOT1_1476 (N4872, N4808);
nand NAND2_1477 (N4873, N4664, N4830);
or OR3_1478 (N4876, N4794, N4797, N4341);
nor NOR3_1479 (N4880, N4794, N4797, N4341);
not NOT1_1480 (N4885, N4812);
not NOT1_1481 (N4889, N4822);
nand NAND2_1482 (N4895, N4859, N4860);
not NOT1_1483 (N4896, N4844);
nand NAND2_1484 (N4897, N4844, N4706);
not NOT1_1485 (N4898, N4847);
nand NAND2_1486 (N4899, N4847, N4707);
nor NOR2_1487 (N4900, N4868, N4564);
and AND4_1488 (N4901, N4717, N4757, N4823, N4564);
not NOT1_1489 (N4902, N4850);
not NOT1_1490 (N4904, N4854);
nand NAND2_1491 (N4905, N4854, N4872);
nand NAND2_1492 (N4906, N4873, N4829);
and AND2_1493 (N4907, N4818, N2123);
and AND2_1494 (N4913, N4823, N2125);
and AND2_1495 (N4916, N4818, N4644);
not NOT1_1496 (N4920, N4880);
and AND2_1497 (N4921, N4895, N2184);
nand NAND2_1498 (N4924, N4656, N4896);
nand NAND2_1499 (N4925, N4659, N4898);
or OR2_1500 (N4926, N4900, N4901);
nand NAND2_1501 (N4928, N4889, N4870);
not NOT1_1502 (N4929, N4889);
nand NAND2_1503 (N4930, N4808, N4904);
not NOT1_1504 (N4931, N4906);
buf BUFF1_1505 (N4937, N4876);
buf BUFF1_1506 (N4940, N4876);
and AND2_1507 (N4944, N4876, N4920);
nand NAND2_1508 (N4946, N4924, N4897);
nand NAND2_1509 (N4949, N4925, N4899);
nand NAND2_1510 (N4950, N4916, N4902);
not NOT1_1511 (N4951, N4916);
nand NAND2_1512 (N4952, N4805, N4929);
nand NAND2_1513 (N4953, N4930, N4905);
and AND2_1514 (N4954, N4926, N2737);
and AND2_1515 (N4957, N4931, N2741);
or OR3_1516 (N4964, N2764, N2483, N4921);
nor NOR3_1517 (N4965, N2764, N2483, N4921);
not NOT1_1518 (N4968, N4949);
nand NAND2_1519 (N4969, N4850, N4951);
nand NAND2_1520 (N4970, N4952, N4928);
and AND2_1521 (N4973, N4953, N2739);
not NOT1_1522 (N4978, N4937);
not NOT1_1523 (N4979, N4940);
not NOT1_1524 (N4980, N4965);
nor NOR2_1525 (N4981, N4968, N4722);
and AND4_1526 (N4982, N4818, N4743, N4946, N4722);
nand NAND2_1527 (N4983, N4950, N4969);
not NOT1_1528 (N4984, N4970);
and AND2_1529 (N4985, N4946, N2121);
or OR3_1530 (N4988, N4913, N4954, N4344);
nor NOR3_1531 (N4991, N4913, N4954, N4344);
or OR3_1532 (N4996, N4800, N4957, N4347);
nor NOR3_1533 (N4999, N4800, N4957, N4347);
and AND2_1534 (N5002, N4964, N4980);
or OR2_1535 (N5007, N4981, N4982);
and AND2_1536 (N5010, N4983, N2731);
and AND2_1537 (N5013, N4984, N2733);
or OR3_1538 (N5018, N4838, N4973, N4475);
nor NOR3_1539 (N5021, N4838, N4973, N4475);
not NOT1_1540 (N5026, N4991);
not NOT1_1541 (N5029, N4999);
and AND2_1542 (N5030, N5007, N2729);
buf BUFF1_1543 (N5039, N4996);
buf BUFF1_1544 (N5042, N4988);
and AND2_1545 (N5045, N4988, N5026);
not NOT1_1546 (N5046, N5021);
and AND2_1547 (N5047, N4996, N5029);
or OR3_1548 (N5050, N4831, N5010, N4472);
nor NOR3_1549 (N5055, N4831, N5010, N4472);
or OR3_1550 (N5058, N4907, N5013, N4338);
nor NOR3_1551 (N5061, N4907, N5013, N4338);
and AND4_1552 (N5066, N4730, N4999, N5021, N4991);
buf BUFF1_1553 (N5070, N5018);
and AND2_1554 (N5078, N5018, N5046);
or OR3_1555 (N5080, N4985, N5030, N4335);
nor NOR3_1556 (N5085, N4985, N5030, N4335);
nand NAND2_1557 (N5094, N5039, N4885);
not NOT1_1558 (N5095, N5039);
not NOT1_1559 (N5097, N5042);
and AND2_1560 (N5102, N5050, N5050);
not NOT1_1561 (N5103, N5061);
nand NAND2_1562 (N5108, N4812, N5095);
not NOT1_1563 (N5109, N5070);
nand NAND2_1564 (N5110, N5070, N5097);
buf BUFF1_1565 (N5111, N5058);
and AND2_1566 (N5114, N5050, N1461);
buf BUFF1_1567 (N5117, N5050);
and AND2_1568 (N5120, N5080, N5080);
and AND2_1569 (N5121, N5058, N5103);
nand NAND2_1570 (N5122, N5094, N5108);
nand NAND2_1571 (N5125, N5042, N5109);
and AND2_1572 (N5128, N1461, N5080);
and AND4_1573 (N5133, N4880, N5061, N5055, N5085);
and AND3_1574 (N5136, N5055, N5085, N1464);
buf BUFF1_1575 (N5139, N5080);
nand NAND2_1576 (N5145, N5125, N5110);
buf BUFF1_1577 (N5151, N5111);
buf BUFF1_1578 (N5154, N5111);
not NOT1_1579 (N5159, N5117);
buf BUFF1_1580 (N5160, N5114);
buf BUFF1_1581 (N5163, N5114);
and AND2_1582 (N5166, N5066, N5133);
and AND2_1583 (N5173, N5066, N5133);
buf BUFF1_1584 (N5174, N5122);
buf BUFF1_1585 (N5177, N5122);
not NOT1_1586 (N5182, N5139);
nand NAND2_1587 (N5183, N5139, N5159);
buf BUFF1_1588 (N5184, N5128);
buf BUFF1_1589 (N5188, N5128);
not NOT1_1590 (N5192, N5166);
nor NOR2_1591 (N5193, N5136, N5173);
nand NAND2_1592 (N5196, N5151, N4978);
not NOT1_1593 (N5197, N5151);
nand NAND2_1594 (N5198, N5154, N4979);
not NOT1_1595 (N5199, N5154);
not NOT1_1596 (N5201, N5160);
not NOT1_1597 (N5203, N5163);
buf BUFF1_1598 (N5205, N5145);
buf BUFF1_1599 (N5209, N5145);
nand NAND2_1600 (N5212, N5117, N5182);
and AND2_1601 (N5215, N213, N5193);
not NOT1_1602 (N5217, N5174);
not NOT1_1603 (N5219, N5177);
nand NAND2_1604 (N5220, N4937, N5197);
nand NAND2_1605 (N5221, N4940, N5199);
not NOT1_1606 (N5222, N5184);
nand NAND2_1607 (N5223, N5184, N5201);
nand NAND2_1608 (N5224, N5188, N5203);
not NOT1_1609 (N5225, N5188);
nand NAND2_1610 (N5228, N5183, N5212);
not NOT1_1611 (N5231, N5215);
nand NAND2_1612 (N5232, N5205, N5217);
not NOT1_1613 (N5233, N5205);
nand NAND2_1614 (N5234, N5209, N5219);
not NOT1_1615 (N5235, N5209);
nand NAND2_1616 (N5236, N5196, N5220);
nand NAND2_1617 (N5240, N5198, N5221);
nand NAND2_1618 (N5242, N5160, N5222);
nand NAND2_1619 (N5243, N5163, N5225);
nand NAND2_1620 (N5245, N5174, N5233);
nand NAND2_1621 (N5246, N5177, N5235);
not NOT1_1622 (N5250, N5240);
not NOT1_1623 (N5253, N5228);
nand NAND2_1624 (N5254, N5242, N5223);
nand NAND2_1625 (N5257, N5243, N5224);
nand NAND2_1626 (N5258, N5232, N5245);
nand NAND2_1627 (N5261, N5234, N5246);
not NOT1_1628 (N5266, N5257);
buf BUFF1_1629 (N5269, N5236);
and AND3_1630 (N5277, N5236, N5254, N2307);
and AND3_1631 (N5278, N5250, N5254, N2310);
not NOT1_1632 (N5279, N5261);
not NOT1_1633 (N5283, N5269);
nand NAND2_1634 (N5284, N5269, N5253);
and AND3_1635 (N5285, N5236, N5266, N2310);
and AND3_1636 (N5286, N5250, N5266, N2307);
buf BUFF1_1637 (N5289, N5258);
buf BUFF1_1638 (N5292, N5258);
nand NAND2_1639 (N5295, N5228, N5283);
or OR4_1640 (N5298, N5277, N5285, N5278, N5286);
buf BUFF1_1641 (N5303, N5279);
buf BUFF1_1642 (N5306, N5279);
nand NAND2_1643 (N5309, N5295, N5284);
not NOT1_1644 (N5312, N5292);
not NOT1_1645 (N5313, N5289);
not NOT1_1646 (N5322, N5306);
not NOT1_1647 (N5323, N5303);
buf BUFF1_1648 (N5324, N5298);
buf BUFF1_1649 (N5327, N5298);
buf BUFF1_1650 (N5332, N5309);
buf BUFF1_1651 (N5335, N5309);
nand NAND2_1652 (N5340, N5324, N5323);
nand NAND2_1653 (N5341, N5327, N5322);
not NOT1_1654 (N5344, N5327);
not NOT1_1655 (N5345, N5324);
nand NAND2_1656 (N5348, N5332, N5313);
nand NAND2_1657 (N5349, N5335, N5312);
nand NAND2_1658 (N5350, N5303, N5345);
nand NAND2_1659 (N5351, N5306, N5344);
not NOT1_1660 (N5352, N5335);
not NOT1_1661 (N5353, N5332);
nand NAND2_1662 (N5354, N5289, N5353);
nand NAND2_1663 (N5355, N5292, N5352);
nand NAND2_1664 (N5356, N5350, N5340);
nand NAND2_1665 (N5357, N5351, N5341);
nand NAND2_1666 (N5358, N5348, N5354);
nand NAND2_1667 (N5359, N5349, N5355);
and AND2_1668 (N5360, N5356, N5357);
nand NAND2_1669 (N5361, N5358, N5359);

endmodule